<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.28" registration="Bezirksschwimmverband Südwestsachsen">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Marienberg" course="SCM" name="28. Internationaler Erzgebirgs-Schwimmcup 2025" nation="GER" organizer="Schwimm-Team Erzgebirge e.V." hostclub="Schwimm-Team Erzgebirge e.V." deadline="2025-12-02" timing="AUTOMATIC">
      <CONTACT city="Olbernhau" email="alex@schwimmteamerzgebirge.de" internet="www.erzgebirgsschwimmcup.de" name="Steiner, Alexander" phone="+49 373607 5177" street="Hammergasse 24" zip="09526" />
      <AGEDATE type="YEAR" value="2025-01-01" />
      <SESSIONS>
        <SESSION number="1" date="2025-12-13" daytime="08:45" officialmeeting="08:15" warmupfrom="07:30">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="F" round="TIM" order="1">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="1001" number="1" daytime="08:45" />
                <HEAT heatid="1002" number="2" daytime="08:47" />
                <HEAT heatid="1003" number="3" daytime="08:49" />
                <HEAT heatid="1004" number="4" daytime="08:51" />
                <HEAT heatid="1005" number="5" daytime="08:53" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="1" resultid="964" />
                    <RANKING place="2" resultid="1074" />
                    <RANKING place="5" resultid="1391" />
                    <RANKING place="3" resultid="1482" />
                    <RANKING place="4" resultid="1819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="7" resultid="211" />
                    <RANKING place="1" resultid="250" />
                    <RANKING place="8" resultid="503" />
                    <RANKING place="3" resultid="907" />
                    <RANKING place="6" resultid="1026" />
                    <RANKING place="2" resultid="1103" />
                    <RANKING place="5" resultid="1408" />
                    <RANKING place="4" resultid="1772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="1321" />
                    <RANKING place="1" resultid="1476" />
                    <RANKING place="2" resultid="1535" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="2" gender="M" round="TIM" order="2">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="2001" number="1" daytime="08:58" />
                <HEAT heatid="2002" number="2" daytime="09:00" />
                <HEAT heatid="2003" number="3" daytime="09:02" />
                <HEAT heatid="2004" number="4" daytime="09:04" />
                <HEAT heatid="2005" number="5" daytime="09:06" />
                <HEAT heatid="2006" number="6" daytime="09:08" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="1" resultid="996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="7" resultid="285" />
                    <RANKING place="1" resultid="544" />
                    <RANKING place="5" resultid="555" />
                    <RANKING place="2" resultid="1064" />
                    <RANKING place="4" resultid="1140" />
                    <RANKING place="3" resultid="1420" />
                    <RANKING place="6" resultid="1541" />
                    <RANKING place="8" resultid="2216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="6" />
                    <RANKING place="3" resultid="113" />
                    <RANKING place="1" resultid="437" />
                    <RANKING place="4" resultid="1218" />
                    <RANKING place="6" resultid="2011" />
                    <RANKING place="7" resultid="2046" />
                    <RANKING place="5" resultid="2152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="262" />
                    <RANKING place="5" resultid="722" />
                    <RANKING place="1" resultid="800" />
                    <RANKING place="4" resultid="1208" />
                    <RANKING place="2" resultid="1278" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="3" gender="F" round="TIM" order="3">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="3000" number="0" />
                <HEAT heatid="3001" number="1" daytime="09:13" />
                <HEAT heatid="3002" number="2" daytime="09:15" />
                <HEAT heatid="3003" number="3" daytime="09:16" />
                <HEAT heatid="3004" number="4" daytime="09:17" />
                <HEAT heatid="3005" number="5" daytime="09:19" />
                <HEAT heatid="3006" number="6" daytime="09:20" />
                <HEAT heatid="3007" number="7" daytime="09:21" />
                <HEAT heatid="3008" number="8" daytime="09:23" />
                <HEAT heatid="3009" number="9" daytime="09:24" />
                <HEAT heatid="3010" number="10" daytime="09:25" />
                <HEAT heatid="3011" number="11" daytime="09:26" />
                <HEAT heatid="3012" number="12" daytime="09:28" />
                <HEAT heatid="3013" number="13" daytime="09:29" />
                <HEAT heatid="3014" number="14" daytime="09:30" />
                <HEAT heatid="3015" number="15" daytime="09:31" />
                <HEAT heatid="3016" number="16" daytime="09:32" />
                <HEAT heatid="3017" number="17" daytime="09:33" />
                <HEAT heatid="3018" number="18" daytime="09:34" />
                <HEAT heatid="3019" number="19" daytime="09:35" />
                <HEAT heatid="3020" number="20" daytime="09:37" />
                <HEAT heatid="3021" number="21" daytime="09:38" />
                <HEAT heatid="3022" number="22" daytime="09:39" />
                <HEAT heatid="3023" number="23" daytime="09:40" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="12" resultid="312" />
                    <RANKING place="14" resultid="393" />
                    <RANKING place="7" resultid="451" />
                    <RANKING place="17" resultid="690" />
                    <RANKING place="13" resultid="863" />
                    <RANKING place="5" resultid="876" />
                    <RANKING place="1" resultid="894" />
                    <RANKING place="11" resultid="922" />
                    <RANKING place="16" resultid="1084" />
                    <RANKING place="2" resultid="1295" />
                    <RANKING place="9" resultid="1369" />
                    <RANKING place="4" resultid="1494" />
                    <RANKING place="3" resultid="1551" />
                    <RANKING place="6" resultid="1712" />
                    <RANKING place="15" resultid="1897" />
                    <RANKING place="8" resultid="1941" />
                    <RANKING place="10" resultid="1969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="9" resultid="11" />
                    <RANKING place="10" resultid="36" />
                    <RANKING place="3" resultid="40" />
                    <RANKING place="11" resultid="45" />
                    <RANKING place="15" resultid="239" />
                    <RANKING place="2" resultid="353" />
                    <RANKING place="5" resultid="590" />
                    <RANKING place="7" resultid="696" />
                    <RANKING place="1" resultid="867" />
                    <RANKING place="19" resultid="880" />
                    <RANKING place="16" resultid="884" />
                    <RANKING place="20" resultid="898" />
                    <RANKING place="13" resultid="1002" />
                    <RANKING place="6" resultid="1289" />
                    <RANKING place="8" resultid="1426" />
                    <RANKING place="12" resultid="1444" />
                    <RANKING place="14" resultid="1516" />
                    <RANKING place="17" resultid="1835" />
                    <RANKING place="18" resultid="2105" />
                    <RANKING place="4" resultid="2117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="205" />
                    <RANKING place="1" resultid="298" />
                    <RANKING place="9" resultid="317" />
                    <RANKING place="7" resultid="716" />
                    <RANKING place="17" resultid="871" />
                    <RANKING place="14" resultid="1050" />
                    <RANKING place="8" resultid="1075" />
                    <RANKING place="6" resultid="1162" />
                    <RANKING place="10" resultid="1315" />
                    <RANKING place="5" resultid="1373" />
                    <RANKING place="4" resultid="1483" />
                    <RANKING place="12" resultid="1510" />
                    <RANKING place="2" resultid="1651" />
                    <RANKING place="11" resultid="1657" />
                    <RANKING place="13" resultid="2025" />
                    <RANKING place="15" resultid="2140" />
                    <RANKING place="16" resultid="2188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="4" resultid="193" />
                    <RANKING place="3" resultid="199" />
                    <RANKING place="5" resultid="888" />
                    <RANKING place="6" resultid="1010" />
                    <RANKING place="8" resultid="1021" />
                    <RANKING place="1" resultid="1488" />
                    <RANKING place="7" resultid="1546" />
                    <RANKING place="2" resultid="1773" />
                    <RANKING place="11" resultid="1987" />
                    <RANKING place="10" resultid="2130" />
                    <RANKING place="9" resultid="2135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="13" resultid="187" />
                    <RANKING place="5" resultid="244" />
                    <RANKING place="1" resultid="457" />
                    <RANKING place="2" resultid="672" />
                    <RANKING place="6" resultid="728" />
                    <RANKING place="15" resultid="980" />
                    <RANKING place="12" resultid="1169" />
                    <RANKING place="10" resultid="1183" />
                    <RANKING place="4" resultid="1228" />
                    <RANKING place="11" resultid="1385" />
                    <RANKING place="8" resultid="1466" />
                    <RANKING place="3" resultid="1536" />
                    <RANKING place="18" resultid="1568" />
                    <RANKING place="16" resultid="1883" />
                    <RANKING place="17" resultid="1963" />
                    <RANKING place="14" resultid="2004" />
                    <RANKING place="7" resultid="2123" />
                    <RANKING place="9" resultid="2229" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="4" gender="M" round="TIM" order="4">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="4000" number="0" />
                <HEAT heatid="4001" number="1" daytime="09:44" />
                <HEAT heatid="4002" number="2" daytime="09:45" />
                <HEAT heatid="4003" number="3" daytime="09:47" />
                <HEAT heatid="4004" number="4" daytime="09:48" />
                <HEAT heatid="4005" number="5" daytime="09:49" />
                <HEAT heatid="4006" number="6" daytime="09:51" />
                <HEAT heatid="4007" number="7" daytime="09:52" />
                <HEAT heatid="4008" number="8" daytime="09:53" />
                <HEAT heatid="4009" number="9" daytime="09:54" />
                <HEAT heatid="4010" number="10" daytime="09:55" />
                <HEAT heatid="4011" number="11" daytime="09:56" />
                <HEAT heatid="4012" number="12" daytime="09:58" />
                <HEAT heatid="4013" number="13" daytime="09:59" />
                <HEAT heatid="4014" number="14" daytime="10:00" />
                <HEAT heatid="4015" number="15" daytime="10:01" />
                <HEAT heatid="4016" number="16" daytime="10:02" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="5" resultid="372" />
                    <RANKING place="1" resultid="468" />
                    <RANKING place="4" resultid="481" />
                    <RANKING place="2" resultid="525" />
                    <RANKING place="6" resultid="1056" />
                    <RANKING place="3" resultid="1916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="3" resultid="1" />
                    <RANKING place="8" resultid="20" />
                    <RANKING place="6" resultid="32" />
                    <RANKING place="10" resultid="217" />
                    <RANKING place="1" resultid="322" />
                    <RANKING place="5" resultid="366" />
                    <RANKING place="4" resultid="586" />
                    <RANKING place="9" resultid="734" />
                    <RANKING place="7" resultid="926" />
                    <RANKING place="2" resultid="1645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="6" resultid="228" />
                    <RANKING place="3" resultid="292" />
                    <RANKING place="2" resultid="417" />
                    <RANKING place="1" resultid="668" />
                    <RANKING place="4" resultid="684" />
                    <RANKING place="5" resultid="1525" />
                    <RANKING place="7" resultid="1556" />
                    <RANKING place="8" resultid="2159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="4" resultid="286" />
                    <RANKING place="3" resultid="549" />
                    <RANKING place="5" resultid="556" />
                    <RANKING place="2" resultid="934" />
                    <RANKING place="7" resultid="1141" />
                    <RANKING place="1" resultid="1421" />
                    <RANKING place="6" resultid="1693" />
                    <RANKING place="10" resultid="1716" />
                    <RANKING place="9" resultid="1829" />
                    <RANKING place="8" resultid="1926" />
                    <RANKING place="11" resultid="1999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="181" />
                    <RANKING place="7" resultid="508" />
                    <RANKING place="10" resultid="1080" />
                    <RANKING place="2" resultid="1438" />
                    <RANKING place="11" resultid="1583" />
                    <RANKING place="6" resultid="1602" />
                    <RANKING place="8" resultid="1908" />
                    <RANKING place="5" resultid="2039" />
                    <RANKING place="9" resultid="2047" />
                    <RANKING place="1" resultid="2063" />
                    <RANKING place="4" resultid="2153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="91" />
                    <RANKING place="2" resultid="598" />
                    <RANKING place="5" resultid="602" />
                    <RANKING place="4" resultid="1564" />
                    <RANKING place="3" resultid="1868" />
                    <RANKING place="6" resultid="1921" />
                    <RANKING place="7" resultid="1953" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="5" gender="F" round="TIM" order="5">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="5000" number="0" />
                <HEAT heatid="5001" number="1" daytime="10:06" />
                <HEAT heatid="5002" number="2" daytime="10:09" />
                <HEAT heatid="5003" number="3" daytime="10:12" />
                <HEAT heatid="5004" number="4" daytime="10:14" />
                <HEAT heatid="5005" number="5" daytime="10:17" />
                <HEAT heatid="5006" number="6" daytime="10:19" />
                <HEAT heatid="5007" number="7" daytime="10:21" />
                <HEAT heatid="5008" number="8" daytime="10:23" />
                <HEAT heatid="5009" number="9" daytime="10:25" />
                <HEAT heatid="5010" number="10" daytime="10:27" />
                <HEAT heatid="5011" number="11" daytime="10:29" />
                <HEAT heatid="5012" number="12" daytime="10:32" />
                <HEAT heatid="5013" number="13" daytime="10:34" />
                <HEAT heatid="5014" number="14" daytime="10:36" />
                <HEAT heatid="5015" number="15" daytime="10:38" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="6" resultid="313" />
                    <RANKING place="3" resultid="913" />
                    <RANKING place="1" resultid="1337" />
                    <RANKING place="4" resultid="1530" />
                    <RANKING place="5" resultid="1713" />
                    <RANKING place="7" resultid="1970" />
                    <RANKING place="2" resultid="2257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="7" resultid="24" />
                    <RANKING place="2" resultid="37" />
                    <RANKING place="4" resultid="48" />
                    <RANKING place="8" resultid="562" />
                    <RANKING place="5" resultid="591" />
                    <RANKING place="3" resultid="1173" />
                    <RANKING place="6" resultid="1445" />
                    <RANKING place="1" resultid="1702" />
                    <RANKING place="9" resultid="2059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="4" resultid="299" />
                    <RANKING place="2" resultid="341" />
                    <RANKING place="6" resultid="717" />
                    <RANKING place="9" resultid="872" />
                    <RANKING place="7" resultid="1051" />
                    <RANKING place="3" resultid="1088" />
                    <RANKING place="1" resultid="1300" />
                    <RANKING place="8" resultid="1460" />
                    <RANKING place="5" resultid="1675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="9" resultid="78" />
                    <RANKING place="7" resultid="95" />
                    <RANKING place="2" resultid="109" />
                    <RANKING place="6" resultid="116" />
                    <RANKING place="1" resultid="251" />
                    <RANKING place="4" resultid="347" />
                    <RANKING place="12" resultid="504" />
                    <RANKING place="13" resultid="889" />
                    <RANKING place="8" resultid="908" />
                    <RANKING place="14" resultid="1011" />
                    <RANKING place="16" resultid="1022" />
                    <RANKING place="5" resultid="1027" />
                    <RANKING place="10" resultid="1331" />
                    <RANKING place="3" resultid="1409" />
                    <RANKING place="10" resultid="1432" />
                    <RANKING place="15" resultid="2131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="7" resultid="102" />
                    <RANKING place="6" resultid="188" />
                    <RANKING place="2" resultid="245" />
                    <RANKING place="8" resultid="519" />
                    <RANKING place="10" resultid="729" />
                    <RANKING place="9" resultid="981" />
                    <RANKING place="4" resultid="1184" />
                    <RANKING place="3" resultid="1306" />
                    <RANKING place="1" resultid="1477" />
                    <RANKING place="5" resultid="1884" />
                    <RANKING place="13" resultid="1964" />
                    <RANKING place="12" resultid="2005" />
                    <RANKING place="11" resultid="2224" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="6" gender="M" round="TIM" order="6">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="6000" number="0" />
                <HEAT heatid="6001" number="1" daytime="10:43" />
                <HEAT heatid="6002" number="2" daytime="10:46" />
                <HEAT heatid="6003" number="3" daytime="10:48" />
                <HEAT heatid="6004" number="4" daytime="10:50" />
                <HEAT heatid="6005" number="5" daytime="10:53" />
                <HEAT heatid="6006" number="6" daytime="10:55" />
                <HEAT heatid="6007" number="7" daytime="10:57" />
                <HEAT heatid="6008" number="8" daytime="10:59" />
                <HEAT heatid="6009" number="9" daytime="11:02" />
                <HEAT heatid="6010" number="10" daytime="11:04" />
                <HEAT heatid="6011" number="11" daytime="11:06" />
                <HEAT heatid="6012" number="12" daytime="11:08" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="2" resultid="469" />
                    <RANKING place="4" resultid="482" />
                    <RANKING place="1" resultid="1310" />
                    <RANKING place="3" resultid="1917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="2" resultid="33" />
                    <RANKING place="4" resultid="367" />
                    <RANKING place="5" resultid="752" />
                    <RANKING place="3" resultid="1753" />
                    <RANKING place="1" resultid="1981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="4" resultid="293" />
                    <RANKING place="3" resultid="529" />
                    <RANKING place="6" resultid="685" />
                    <RANKING place="2" resultid="1792" />
                    <RANKING place="5" resultid="2160" />
                    <RANKING place="1" resultid="2250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="3" resultid="404" />
                    <RANKING place="4" resultid="935" />
                    <RANKING place="1" resultid="958" />
                    <RANKING place="2" resultid="990" />
                    <RANKING place="5" resultid="2217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="74" />
                    <RANKING place="1" resultid="438" />
                    <RANKING place="5" resultid="509" />
                    <RANKING place="6" resultid="1909" />
                    <RANKING place="2" resultid="2012" />
                    <RANKING place="3" resultid="2040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="9" resultid="723" />
                    <RANKING place="1" resultid="801" />
                    <RANKING place="5" resultid="1279" />
                    <RANKING place="2" resultid="1397" />
                    <RANKING place="10" resultid="1619" />
                    <RANKING place="6" resultid="1728" />
                    <RANKING place="3" resultid="1814" />
                    <RANKING place="8" resultid="1922" />
                    <RANKING place="7" resultid="1954" />
                    <RANKING place="4" resultid="2279" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="7" gender="F" round="TIM" order="7">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="7000" number="0" />
                <HEAT heatid="7001" number="1" daytime="11:13" />
                <HEAT heatid="7002" number="2" daytime="11:14" />
                <HEAT heatid="7003" number="3" daytime="11:16" />
                <HEAT heatid="7004" number="4" daytime="11:17" />
                <HEAT heatid="7005" number="5" daytime="11:18" />
                <HEAT heatid="7006" number="6" daytime="11:20" />
                <HEAT heatid="7007" number="7" daytime="11:21" />
                <HEAT heatid="7008" number="8" daytime="11:22" />
                <HEAT heatid="7009" number="9" daytime="11:23" />
                <HEAT heatid="7010" number="10" daytime="11:24" />
                <HEAT heatid="7011" number="11" daytime="11:25" />
                <HEAT heatid="7012" number="12" daytime="11:27" />
                <HEAT heatid="7013" number="13" daytime="11:28" />
                <HEAT heatid="7014" number="14" daytime="11:29" />
                <HEAT heatid="7015" number="15" daytime="11:30" />
                <HEAT heatid="7016" number="16" daytime="11:31" />
                <HEAT heatid="7017" number="17" daytime="11:32" />
                <HEAT heatid="7018" number="18" daytime="11:33" />
                <HEAT heatid="7019" number="19" daytime="11:34" />
                <HEAT heatid="7020" number="20" daytime="11:35" />
                <HEAT heatid="7021" number="21" daytime="11:36" />
                <HEAT heatid="7022" number="22" daytime="11:37" />
                <HEAT heatid="7023" number="23" daytime="11:38" />
                <HEAT heatid="7024" number="24" daytime="11:39" />
                <HEAT heatid="7025" number="25" daytime="11:40" />
                <HEAT heatid="7026" number="26" daytime="11:41" />
                <HEAT heatid="7027" number="27" daytime="11:42" />
                <HEAT heatid="7028" number="28" daytime="11:43" />
                <HEAT heatid="7029" number="29" daytime="11:44" />
                <HEAT heatid="7030" number="30" daytime="11:45" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="9" resultid="314" />
                    <RANKING place="15" resultid="394" />
                    <RANKING place="6" resultid="452" />
                    <RANKING place="12" resultid="692" />
                    <RANKING place="10" resultid="864" />
                    <RANKING place="2" resultid="877" />
                    <RANKING place="1" resultid="895" />
                    <RANKING place="16" resultid="923" />
                    <RANKING place="19" resultid="1085" />
                    <RANKING place="7" resultid="1171" />
                    <RANKING place="5" resultid="1296" />
                    <RANKING place="8" resultid="1338" />
                    <RANKING place="13" resultid="1370" />
                    <RANKING place="3" resultid="1495" />
                    <RANKING place="4" resultid="1552" />
                    <RANKING place="11" resultid="1898" />
                    <RANKING place="18" resultid="1942" />
                    <RANKING place="17" resultid="1971" />
                    <RANKING place="14" resultid="2258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="6" resultid="12" />
                    <RANKING place="4" resultid="15" />
                    <RANKING place="18" resultid="25" />
                    <RANKING place="17" resultid="38" />
                    <RANKING place="1" resultid="41" />
                    <RANKING place="19" resultid="46" />
                    <RANKING place="13" resultid="49" />
                    <RANKING place="16" resultid="240" />
                    <RANKING place="3" resultid="354" />
                    <RANKING place="5" resultid="499" />
                    <RANKING place="15" resultid="563" />
                    <RANKING place="7" resultid="697" />
                    <RANKING place="2" resultid="868" />
                    <RANKING place="27" resultid="881" />
                    <RANKING place="26" resultid="885" />
                    <RANKING place="25" resultid="899" />
                    <RANKING place="11" resultid="1174" />
                    <RANKING place="10" resultid="1290" />
                    <RANKING place="9" resultid="1427" />
                    <RANKING place="21" resultid="1446" />
                    <RANKING place="24" resultid="1517" />
                    <RANKING place="12" resultid="1703" />
                    <RANKING place="22" resultid="1778" />
                    <RANKING place="14" resultid="1836" />
                    <RANKING place="23" resultid="2060" />
                    <RANKING place="20" resultid="2106" />
                    <RANKING place="8" resultid="2118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="6" resultid="206" />
                    <RANKING place="8" resultid="300" />
                    <RANKING place="19" resultid="318" />
                    <RANKING place="3" resultid="342" />
                    <RANKING place="14" resultid="595" />
                    <RANKING place="9" resultid="718" />
                    <RANKING place="24" resultid="873" />
                    <RANKING place="10" resultid="965" />
                    <RANKING place="13" resultid="1052" />
                    <RANKING place="12" resultid="1089" />
                    <RANKING place="7" resultid="1163" />
                    <RANKING place="1" resultid="1301" />
                    <RANKING place="18" resultid="1316" />
                    <RANKING place="15" resultid="1374" />
                    <RANKING place="20" resultid="1392" />
                    <RANKING place="21" resultid="1461" />
                    <RANKING place="5" resultid="1484" />
                    <RANKING place="17" resultid="1511" />
                    <RANKING place="4" resultid="1652" />
                    <RANKING place="16" resultid="1658" />
                    <RANKING place="2" resultid="1676" />
                    <RANKING place="11" resultid="1820" />
                    <RANKING place="22" resultid="2026" />
                    <RANKING place="23" resultid="2141" />
                    <RANKING place="25" resultid="2189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="6" resultid="117" />
                    <RANKING place="5" resultid="194" />
                    <RANKING place="7" resultid="200" />
                    <RANKING place="10" resultid="212" />
                    <RANKING place="1" resultid="252" />
                    <RANKING place="9" resultid="348" />
                    <RANKING place="8" resultid="432" />
                    <RANKING place="12" resultid="890" />
                    <RANKING place="15" resultid="1012" />
                    <RANKING place="17" resultid="1023" />
                    <RANKING place="3" resultid="1104" />
                    <RANKING place="13" resultid="1332" />
                    <RANKING place="11" resultid="1433" />
                    <RANKING place="4" resultid="1489" />
                    <RANKING place="14" resultid="1547" />
                    <RANKING place="2" resultid="1774" />
                    <RANKING place="18" resultid="1988" />
                    <RANKING place="19" resultid="2132" />
                    <RANKING place="16" resultid="2136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="11" resultid="103" />
                    <RANKING place="13" resultid="189" />
                    <RANKING place="1" resultid="458" />
                    <RANKING place="3" resultid="673" />
                    <RANKING place="5" resultid="730" />
                    <RANKING place="15" resultid="982" />
                    <RANKING place="6" resultid="1229" />
                    <RANKING place="9" resultid="1307" />
                    <RANKING place="4" resultid="1322" />
                    <RANKING place="12" resultid="1386" />
                    <RANKING place="7" resultid="1467" />
                    <RANKING place="2" resultid="1537" />
                    <RANKING place="16" resultid="1569" />
                    <RANKING place="18" resultid="1965" />
                    <RANKING place="10" resultid="2006" />
                    <RANKING place="8" resultid="2124" />
                    <RANKING place="17" resultid="2225" />
                    <RANKING place="14" resultid="2230" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="8" gender="M" round="TIM" order="8">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="8000" number="0" />
                <HEAT heatid="8001" number="1" daytime="11:49" />
                <HEAT heatid="8002" number="2" daytime="11:50" />
                <HEAT heatid="8003" number="3" daytime="11:52" />
                <HEAT heatid="8004" number="4" daytime="11:53" />
                <HEAT heatid="8005" number="5" daytime="11:54" />
                <HEAT heatid="8006" number="6" daytime="11:55" />
                <HEAT heatid="8007" number="7" daytime="11:56" />
                <HEAT heatid="8008" number="8" daytime="11:58" />
                <HEAT heatid="8009" number="9" daytime="11:59" />
                <HEAT heatid="8010" number="10" daytime="12:00" />
                <HEAT heatid="8011" number="11" daytime="12:01" />
                <HEAT heatid="8012" number="12" daytime="12:02" />
                <HEAT heatid="8013" number="13" daytime="12:03" />
                <HEAT heatid="8014" number="14" daytime="12:04" />
                <HEAT heatid="8015" number="15" daytime="12:05" />
                <HEAT heatid="8016" number="16" daytime="12:06" />
                <HEAT heatid="8017" number="17" daytime="12:07" />
                <HEAT heatid="8018" number="18" daytime="12:08" />
                <HEAT heatid="8019" number="19" daytime="12:09" />
                <HEAT heatid="8020" number="20" daytime="12:09" />
                <HEAT heatid="8021" number="21" daytime="12:11" />
                <HEAT heatid="8022" number="22" daytime="12:12" />
                <HEAT heatid="8023" number="23" daytime="12:13" />
                <HEAT heatid="8024" number="24" daytime="12:14" />
                <HEAT heatid="8025" number="25" daytime="12:14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="5" resultid="373" />
                    <RANKING place="3" resultid="470" />
                    <RANKING place="4" resultid="483" />
                    <RANKING place="1" resultid="526" />
                    <RANKING place="7" resultid="1057" />
                    <RANKING place="6" resultid="1311" />
                    <RANKING place="8" resultid="1826" />
                    <RANKING place="2" resultid="1918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="4" resultid="2" />
                    <RANKING place="14" resultid="21" />
                    <RANKING place="10" resultid="34" />
                    <RANKING place="11" resultid="218" />
                    <RANKING place="2" resultid="323" />
                    <RANKING place="9" resultid="368" />
                    <RANKING place="1" resultid="566" />
                    <RANKING place="5" resultid="587" />
                    <RANKING place="12" resultid="735" />
                    <RANKING place="15" resultid="753" />
                    <RANKING place="6" resultid="927" />
                    <RANKING place="3" resultid="1646" />
                    <RANKING place="7" resultid="1699" />
                    <RANKING place="13" resultid="1769" />
                    <RANKING place="8" resultid="1982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="8" resultid="229" />
                    <RANKING place="4" resultid="418" />
                    <RANKING place="2" resultid="530" />
                    <RANKING place="7" resultid="686" />
                    <RANKING place="5" resultid="997" />
                    <RANKING place="6" resultid="1526" />
                    <RANKING place="9" resultid="1557" />
                    <RANKING place="3" resultid="1793" />
                    <RANKING place="10" resultid="2161" />
                    <RANKING place="1" resultid="2251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="6" resultid="287" />
                    <RANKING place="12" resultid="405" />
                    <RANKING place="1" resultid="545" />
                    <RANKING place="4" resultid="550" />
                    <RANKING place="8" resultid="936" />
                    <RANKING place="5" resultid="959" />
                    <RANKING place="3" resultid="991" />
                    <RANKING place="2" resultid="1065" />
                    <RANKING place="7" resultid="1422" />
                    <RANKING place="10" resultid="1542" />
                    <RANKING place="20" resultid="1618" />
                    <RANKING place="17" resultid="1623" />
                    <RANKING place="13" resultid="1627" />
                    <RANKING place="16" resultid="1631" />
                    <RANKING place="9" resultid="1694" />
                    <RANKING place="18" resultid="1718" />
                    <RANKING place="11" resultid="1830" />
                    <RANKING place="14" resultid="1927" />
                    <RANKING place="19" resultid="2000" />
                    <RANKING place="15" resultid="2218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="7" resultid="7" />
                    <RANKING place="3" resultid="114" />
                    <RANKING place="5" resultid="182" />
                    <RANKING place="2" resultid="439" />
                    <RANKING place="12" resultid="510" />
                    <RANKING place="16" resultid="1081" />
                    <RANKING place="1" resultid="1219" />
                    <RANKING place="6" resultid="1439" />
                    <RANKING place="15" resultid="1584" />
                    <RANKING place="11" resultid="1603" />
                    <RANKING place="14" resultid="1910" />
                    <RANKING place="9" resultid="2013" />
                    <RANKING place="10" resultid="2041" />
                    <RANKING place="13" resultid="2048" />
                    <RANKING place="4" resultid="2064" />
                    <RANKING place="8" resultid="2154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="11" resultid="92" />
                    <RANKING place="3" resultid="263" />
                    <RANKING place="5" resultid="599" />
                    <RANKING place="9" resultid="603" />
                    <RANKING place="13" resultid="724" />
                    <RANKING place="1" resultid="1209" />
                    <RANKING place="2" resultid="1398" />
                    <RANKING place="14" resultid="1565" />
                    <RANKING place="15" resultid="1615" />
                    <RANKING place="8" resultid="1729" />
                    <RANKING place="4" resultid="1815" />
                    <RANKING place="6" resultid="1870" />
                    <RANKING place="10" resultid="1923" />
                    <RANKING place="12" resultid="1955" />
                    <RANKING place="7" resultid="2280" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="9" gender="F" round="TIM" order="9">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="9000" number="0" />
                <HEAT heatid="9001" number="1" daytime="12:18" />
                <HEAT heatid="9002" number="2" daytime="12:21" />
                <HEAT heatid="9003" number="3" daytime="12:23" />
                <HEAT heatid="9004" number="4" daytime="12:26" />
                <HEAT heatid="9005" number="5" daytime="12:28" />
                <HEAT heatid="9006" number="6" daytime="12:30" />
                <HEAT heatid="9007" number="7" daytime="12:32" />
                <HEAT heatid="9008" number="8" daytime="12:34" />
                <HEAT heatid="9009" number="9" daytime="12:36" />
                <HEAT heatid="9010" number="10" daytime="12:38" />
                <HEAT heatid="9011" number="11" daytime="12:40" />
                <HEAT heatid="9012" number="12" daytime="12:42" />
                <HEAT heatid="9013" number="13" daytime="12:44" />
                <HEAT heatid="9014" number="14" daytime="12:46" />
                <HEAT heatid="9015" number="15" daytime="12:48" />
                <HEAT heatid="9016" number="16" daytime="12:50" />
                <HEAT heatid="9017" number="17" daytime="12:52" />
                <HEAT heatid="9018" number="18" daytime="12:54" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="6" resultid="453" />
                    <RANKING place="3" resultid="914" />
                    <RANKING place="4" resultid="1297" />
                    <RANKING place="2" resultid="1339" />
                    <RANKING place="7" resultid="1371" />
                    <RANKING place="1" resultid="1496" />
                    <RANKING place="8" resultid="1531" />
                    <RANKING place="5" resultid="1553" />
                    <RANKING place="9" resultid="1943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="1" resultid="42" />
                    <RANKING place="4" resultid="355" />
                    <RANKING place="5" resultid="500" />
                    <RANKING place="6" resultid="1291" />
                    <RANKING place="2" resultid="1428" />
                    <RANKING place="9" resultid="1518" />
                    <RANKING place="8" resultid="1779" />
                    <RANKING place="7" resultid="2107" />
                    <RANKING place="3" resultid="2119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="7" resultid="207" />
                    <RANKING place="14" resultid="319" />
                    <RANKING place="5" resultid="343" />
                    <RANKING place="4" resultid="966" />
                    <RANKING place="3" resultid="1076" />
                    <RANKING place="6" resultid="1090" />
                    <RANKING place="1" resultid="1302" />
                    <RANKING place="10" resultid="1317" />
                    <RANKING place="12" resultid="1375" />
                    <RANKING place="11" resultid="1393" />
                    <RANKING place="17" resultid="1462" />
                    <RANKING place="13" resultid="1512" />
                    <RANKING place="2" resultid="1653" />
                    <RANKING place="15" resultid="1659" />
                    <RANKING place="8" resultid="1677" />
                    <RANKING place="9" resultid="1821" />
                    <RANKING place="16" resultid="2027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="13" resultid="79" />
                    <RANKING place="9" resultid="96" />
                    <RANKING place="1" resultid="110" />
                    <RANKING place="10" resultid="195" />
                    <RANKING place="8" resultid="201" />
                    <RANKING place="15" resultid="213" />
                    <RANKING place="11" resultid="349" />
                    <RANKING place="7" resultid="433" />
                    <RANKING place="12" resultid="505" />
                    <RANKING place="3" resultid="909" />
                    <RANKING place="6" resultid="1028" />
                    <RANKING place="2" resultid="1105" />
                    <RANKING place="16" resultid="1333" />
                    <RANKING place="4" resultid="1410" />
                    <RANKING place="14" resultid="1434" />
                    <RANKING place="5" resultid="1490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="7" resultid="246" />
                    <RANKING place="4" resultid="459" />
                    <RANKING place="14" resultid="520" />
                    <RANKING place="3" resultid="674" />
                    <RANKING place="8" resultid="1185" />
                    <RANKING place="5" resultid="1230" />
                    <RANKING place="6" resultid="1323" />
                    <RANKING place="11" resultid="1387" />
                    <RANKING place="9" resultid="1468" />
                    <RANKING place="1" resultid="1478" />
                    <RANKING place="2" resultid="1538" />
                    <RANKING place="15" resultid="1886" />
                    <RANKING place="12" resultid="2007" />
                    <RANKING place="13" resultid="2125" />
                    <RANKING place="10" resultid="2231" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="10" number="10" gender="M" round="TIM" order="10">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="10000" number="0" />
                <HEAT heatid="10001" number="1" daytime="12:59" />
                <HEAT heatid="10002" number="2" daytime="13:01" />
                <HEAT heatid="10003" number="3" daytime="13:03" />
                <HEAT heatid="10004" number="4" daytime="13:05" />
                <HEAT heatid="10005" number="5" daytime="13:07" />
                <HEAT heatid="10006" number="6" daytime="13:09" />
                <HEAT heatid="10007" number="7" daytime="13:11" />
                <HEAT heatid="10008" number="8" daytime="13:13" />
                <HEAT heatid="10009" number="9" daytime="13:15" />
                <HEAT heatid="10010" number="10" daytime="13:18" />
                <HEAT heatid="10011" number="11" daytime="13:19" />
                <HEAT heatid="10012" number="12" daytime="13:21" />
                <HEAT heatid="10013" number="13" daytime="13:23" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="1" resultid="374" />
                    <RANKING place="2" resultid="1312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="6" resultid="219" />
                    <RANKING place="2" resultid="324" />
                    <RANKING place="1" resultid="567" />
                    <RANKING place="3" resultid="1647" />
                    <RANKING place="5" resultid="1754" />
                    <RANKING place="4" resultid="1983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="5" resultid="419" />
                    <RANKING place="2" resultid="531" />
                    <RANKING place="6" resultid="669" />
                    <RANKING place="4" resultid="998" />
                    <RANKING place="7" resultid="1527" />
                    <RANKING place="1" resultid="1794" />
                    <RANKING place="3" resultid="2252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="8" resultid="288" />
                    <RANKING place="9" resultid="406" />
                    <RANKING place="1" resultid="546" />
                    <RANKING place="2" resultid="551" />
                    <RANKING place="7" resultid="557" />
                    <RANKING place="4" resultid="960" />
                    <RANKING place="5" resultid="992" />
                    <RANKING place="3" resultid="1066" />
                    <RANKING place="6" resultid="1142" />
                    <RANKING place="11" resultid="1543" />
                    <RANKING place="10" resultid="1831" />
                    <RANKING place="12" resultid="1928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="8" />
                    <RANKING place="4" resultid="183" />
                    <RANKING place="1" resultid="440" />
                    <RANKING place="2" resultid="1440" />
                    <RANKING place="8" resultid="1911" />
                    <RANKING place="6" resultid="2014" />
                    <RANKING place="9" resultid="2049" />
                    <RANKING place="5" resultid="2065" />
                    <RANKING place="7" resultid="2155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="264" />
                    <RANKING place="2" resultid="1399" />
                    <RANKING place="3" resultid="1816" />
                    <RANKING place="5" resultid="1956" />
                    <RANKING place="4" resultid="2281" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="11" gender="X" round="TIM" order="11">
              <SWIMSTYLE stroke="FREE" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="11000" number="0" />
                <HEAT heatid="11001" number="1" daytime="13:28" />
                <HEAT heatid="11002" number="2" daytime="13:31" />
                <HEAT heatid="11003" number="3" daytime="13:33" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="13" agemin="8" name="Jahrgänge 2012 bis 2017">
                  <RANKINGS>
                    <RANKING place="11" resultid="178" />
                    <RANKING place="3" resultid="179" />
                    <RANKING place="4" resultid="279" />
                    <RANKING place="5" resultid="849" />
                    <RANKING place="10" resultid="855" />
                    <RANKING place="7" resultid="856" />
                    <RANKING place="1" resultid="1182" />
                    <RANKING place="2" resultid="1287" />
                    <RANKING place="6" resultid="1849" />
                    <RANKING place="8" resultid="1855" />
                    <RANKING place="9" resultid="1861" />
                    <RANKING place="12" resultid="1865" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2025-12-13" daytime="00:30">
          <EVENTS>
            <EVENT eventid="13" number="12" gender="F" round="TIM" order="12">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="13000" number="0" />
                <HEAT heatid="13001" number="1" daytime="14:09" />
                <HEAT heatid="13002" number="2" daytime="14:11" />
                <HEAT heatid="13003" number="3" daytime="14:12" />
                <HEAT heatid="13004" number="4" daytime="14:13" />
                <HEAT heatid="13005" number="5" daytime="14:14" />
                <HEAT heatid="13006" number="6" daytime="14:16" />
                <HEAT heatid="13007" number="7" daytime="14:17" />
                <HEAT heatid="13008" number="8" daytime="14:18" />
                <HEAT heatid="13009" number="9" daytime="14:19" />
                <HEAT heatid="13010" number="10" daytime="14:20" />
                <HEAT heatid="13011" number="11" daytime="14:21" />
                <HEAT heatid="13012" number="12" daytime="14:22" />
                <HEAT heatid="13013" number="13" daytime="14:24" />
                <HEAT heatid="13014" number="14" daytime="14:25" />
                <HEAT heatid="13015" number="15" daytime="14:26" />
                <HEAT heatid="13016" number="16" daytime="14:27" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="6" resultid="454" />
                    <RANKING place="4" resultid="915" />
                    <RANKING place="2" resultid="1298" />
                    <RANKING place="3" resultid="1340" />
                    <RANKING place="5" resultid="1372" />
                    <RANKING place="1" resultid="1497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="2" resultid="16" />
                    <RANKING place="4" resultid="43" />
                    <RANKING place="7" resultid="50" />
                    <RANKING place="8" resultid="356" />
                    <RANKING place="9" resultid="501" />
                    <RANKING place="6" resultid="564" />
                    <RANKING place="5" resultid="699" />
                    <RANKING place="1" resultid="869" />
                    <RANKING place="10" resultid="1292" />
                    <RANKING place="3" resultid="1429" />
                    <RANKING place="11" resultid="2108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="5" resultid="208" />
                    <RANKING place="9" resultid="320" />
                    <RANKING place="2" resultid="344" />
                    <RANKING place="6" resultid="596" />
                    <RANKING place="4" resultid="967" />
                    <RANKING place="1" resultid="1077" />
                    <RANKING place="8" resultid="1164" />
                    <RANKING place="11" resultid="1394" />
                    <RANKING place="10" resultid="1463" />
                    <RANKING place="3" resultid="1485" />
                    <RANKING place="13" resultid="1513" />
                    <RANKING place="12" resultid="1660" />
                    <RANKING place="7" resultid="1822" />
                    <RANKING place="14" resultid="2028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="7" resultid="196" />
                    <RANKING place="6" resultid="202" />
                    <RANKING place="12" resultid="214" />
                    <RANKING place="1" resultid="253" />
                    <RANKING place="9" resultid="434" />
                    <RANKING place="2" resultid="910" />
                    <RANKING place="3" resultid="1106" />
                    <RANKING place="13" resultid="1334" />
                    <RANKING place="5" resultid="1411" />
                    <RANKING place="10" resultid="1435" />
                    <RANKING place="8" resultid="1491" />
                    <RANKING place="11" resultid="1548" />
                    <RANKING place="4" resultid="1775" />
                    <RANKING place="14" resultid="2137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="9" resultid="190" />
                    <RANKING place="7" resultid="247" />
                    <RANKING place="5" resultid="460" />
                    <RANKING place="12" resultid="521" />
                    <RANKING place="3" resultid="675" />
                    <RANKING place="13" resultid="983" />
                    <RANKING place="6" resultid="1186" />
                    <RANKING place="4" resultid="1324" />
                    <RANKING place="8" resultid="1388" />
                    <RANKING place="1" resultid="1479" />
                    <RANKING place="2" resultid="1539" />
                    <RANKING place="14" resultid="1966" />
                    <RANKING place="11" resultid="2008" />
                    <RANKING place="10" resultid="2232" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="14" number="13" gender="M" round="TIM" order="13">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="14001" number="1" daytime="14:31" />
                <HEAT heatid="14002" number="2" daytime="14:32" />
                <HEAT heatid="14003" number="3" daytime="14:34" />
                <HEAT heatid="14004" number="4" daytime="14:35" />
                <HEAT heatid="14005" number="5" daytime="14:36" />
                <HEAT heatid="14006" number="6" daytime="14:37" />
                <HEAT heatid="14007" number="7" daytime="14:38" />
                <HEAT heatid="14008" number="8" daytime="14:39" />
                <HEAT heatid="14009" number="9" daytime="14:41" />
                <HEAT heatid="14010" number="10" daytime="14:42" />
                <HEAT heatid="14011" number="11" daytime="14:43" />
                <HEAT heatid="14012" number="12" daytime="14:44" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017" />
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="4" resultid="3" />
                    <RANKING place="2" resultid="325" />
                    <RANKING place="5" resultid="369" />
                    <RANKING place="1" resultid="568" />
                    <RANKING place="7" resultid="928" />
                    <RANKING place="3" resultid="1648" />
                    <RANKING place="6" resultid="1984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="4" resultid="420" />
                    <RANKING place="3" resultid="532" />
                    <RANKING place="2" resultid="999" />
                    <RANKING place="1" resultid="2253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="9" resultid="289" />
                    <RANKING place="8" resultid="407" />
                    <RANKING place="1" resultid="547" />
                    <RANKING place="3" resultid="552" />
                    <RANKING place="7" resultid="558" />
                    <RANKING place="12" resultid="937" />
                    <RANKING place="6" resultid="993" />
                    <RANKING place="2" resultid="1067" />
                    <RANKING place="5" resultid="1143" />
                    <RANKING place="4" resultid="1423" />
                    <RANKING place="9" resultid="1544" />
                    <RANKING place="11" resultid="1929" />
                    <RANKING place="14" resultid="2001" />
                    <RANKING place="13" resultid="2219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="9" />
                    <RANKING place="6" resultid="184" />
                    <RANKING place="1" resultid="441" />
                    <RANKING place="2" resultid="1220" />
                    <RANKING place="8" resultid="1441" />
                    <RANKING place="9" resultid="2015" />
                    <RANKING place="7" resultid="2042" />
                    <RANKING place="10" resultid="2050" />
                    <RANKING place="4" resultid="2066" />
                    <RANKING place="5" resultid="2156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="265" />
                    <RANKING place="3" resultid="1210" />
                    <RANKING place="1" resultid="1280" />
                    <RANKING place="2" resultid="1400" />
                    <RANKING place="5" resultid="1957" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="15" number="14" gender="F" round="TIM" order="14">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="15000" number="0" />
                <HEAT heatid="15001" number="1" daytime="14:48" />
                <HEAT heatid="15002" number="2" daytime="14:51" />
                <HEAT heatid="15003" number="3" daytime="14:53" />
                <HEAT heatid="15004" number="4" daytime="14:56" />
                <HEAT heatid="15005" number="5" daytime="14:59" />
                <HEAT heatid="15006" number="6" daytime="15:01" />
                <HEAT heatid="15007" number="7" daytime="15:03" />
                <HEAT heatid="15008" number="8" daytime="15:05" />
                <HEAT heatid="15009" number="9" daytime="15:08" />
                <HEAT heatid="15010" number="10" daytime="15:10" />
                <HEAT heatid="15011" number="11" daytime="15:12" />
                <HEAT heatid="15012" number="12" daytime="15:14" />
                <HEAT heatid="15013" number="13" daytime="15:16" />
                <HEAT heatid="15014" number="14" daytime="15:17" />
                <HEAT heatid="15015" number="15" daytime="15:19" />
                <HEAT heatid="15016" number="16" daytime="15:22" />
                <HEAT heatid="15017" number="17" daytime="15:24" />
                <HEAT heatid="15018" number="18" daytime="15:26" />
                <HEAT heatid="15019" number="19" daytime="15:27" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="9" resultid="395" />
                    <RANKING place="4" resultid="455" />
                    <RANKING place="7" resultid="693" />
                    <RANKING place="11" resultid="1086" />
                    <RANKING place="2" resultid="1299" />
                    <RANKING place="1" resultid="1498" />
                    <RANKING place="5" resultid="1532" />
                    <RANKING place="3" resultid="1554" />
                    <RANKING place="10" resultid="1899" />
                    <RANKING place="8" resultid="1944" />
                    <RANKING place="6" resultid="1972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="7" resultid="13" />
                    <RANKING place="2" resultid="17" />
                    <RANKING place="10" resultid="241" />
                    <RANKING place="1" resultid="357" />
                    <RANKING place="3" resultid="592" />
                    <RANKING place="6" resultid="700" />
                    <RANKING place="4" resultid="1293" />
                    <RANKING place="8" resultid="1519" />
                    <RANKING place="9" resultid="1837" />
                    <RANKING place="11" resultid="2109" />
                    <RANKING place="5" resultid="2120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="4" resultid="209" />
                    <RANKING place="1" resultid="301" />
                    <RANKING place="10" resultid="321" />
                    <RANKING place="9" resultid="597" />
                    <RANKING place="7" resultid="719" />
                    <RANKING place="16" resultid="874" />
                    <RANKING place="3" resultid="968" />
                    <RANKING place="11" resultid="1053" />
                    <RANKING place="2" resultid="1303" />
                    <RANKING place="8" resultid="1318" />
                    <RANKING place="6" resultid="1376" />
                    <RANKING place="13" resultid="1395" />
                    <RANKING place="5" resultid="1486" />
                    <RANKING place="12" resultid="1514" />
                    <RANKING place="15" resultid="1661" />
                    <RANKING place="14" resultid="2029" />
                    <RANKING place="17" resultid="2142" />
                    <RANKING place="18" resultid="2190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="7" resultid="197" />
                    <RANKING place="6" resultid="203" />
                    <RANKING place="1" resultid="254" />
                    <RANKING place="8" resultid="506" />
                    <RANKING place="9" resultid="891" />
                    <RANKING place="5" resultid="911" />
                    <RANKING place="10" resultid="1013" />
                    <RANKING place="12" resultid="1024" />
                    <RANKING place="2" resultid="1107" />
                    <RANKING place="3" resultid="1492" />
                    <RANKING place="11" resultid="1549" />
                    <RANKING place="4" resultid="1776" />
                    <RANKING place="14" resultid="2133" />
                    <RANKING place="13" resultid="2138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="8" resultid="248" />
                    <RANKING place="1" resultid="461" />
                    <RANKING place="7" resultid="731" />
                    <RANKING place="3" resultid="1231" />
                    <RANKING place="4" resultid="1308" />
                    <RANKING place="5" resultid="1325" />
                    <RANKING place="11" resultid="1389" />
                    <RANKING place="6" resultid="1469" />
                    <RANKING place="2" resultid="1540" />
                    <RANKING place="10" resultid="2126" />
                    <RANKING place="12" resultid="2226" />
                    <RANKING place="9" resultid="2233" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="16" number="15" gender="M" round="TIM" order="15">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="16000" number="0" />
                <HEAT heatid="16001" number="1" daytime="15:32" />
                <HEAT heatid="16002" number="2" daytime="15:35" />
                <HEAT heatid="16003" number="3" daytime="15:37" />
                <HEAT heatid="16004" number="4" daytime="15:39" />
                <HEAT heatid="16005" number="5" daytime="15:41" />
                <HEAT heatid="16006" number="6" daytime="15:43" />
                <HEAT heatid="16007" number="7" daytime="15:46" />
                <HEAT heatid="16008" number="8" daytime="15:48" />
                <HEAT heatid="16009" number="9" daytime="15:50" />
                <HEAT heatid="16010" number="10" daytime="15:52" />
                <HEAT heatid="16011" number="11" daytime="15:54" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="3" resultid="375" />
                    <RANKING place="1" resultid="471" />
                    <RANKING place="2" resultid="484" />
                    <RANKING place="4" resultid="1827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="2" resultid="4" />
                    <RANKING place="4" resultid="326" />
                    <RANKING place="1" resultid="569" />
                    <RANKING place="3" resultid="1649" />
                    <RANKING place="5" resultid="1770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="5" resultid="231" />
                    <RANKING place="2" resultid="295" />
                    <RANKING place="1" resultid="421" />
                    <RANKING place="3" resultid="687" />
                    <RANKING place="4" resultid="1528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="4" resultid="408" />
                    <RANKING place="3" resultid="559" />
                    <RANKING place="2" resultid="938" />
                    <RANKING place="5" resultid="1144" />
                    <RANKING place="1" resultid="1424" />
                    <RANKING place="6" resultid="1696" />
                    <RANKING place="9" resultid="1719" />
                    <RANKING place="7" resultid="1832" />
                    <RANKING place="8" resultid="1930" />
                    <RANKING place="10" resultid="2002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="75" />
                    <RANKING place="1" resultid="185" />
                    <RANKING place="4" resultid="1082" />
                    <RANKING place="2" resultid="2067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="93" />
                    <RANKING place="3" resultid="600" />
                    <RANKING place="4" resultid="604" />
                    <RANKING place="6" resultid="725" />
                    <RANKING place="5" resultid="1871" />
                    <RANKING place="1" resultid="2282" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="17" number="16" gender="F" round="TIM" order="16">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="17000" number="0" />
                <HEAT heatid="17001" number="1" daytime="15:59" />
                <HEAT heatid="17002" number="2" daytime="16:00" />
                <HEAT heatid="17003" number="3" daytime="16:02" />
                <HEAT heatid="17004" number="4" daytime="16:04" />
                <HEAT heatid="17005" number="5" daytime="16:05" />
                <HEAT heatid="17006" number="6" daytime="16:06" />
                <HEAT heatid="17007" number="7" daytime="16:08" />
                <HEAT heatid="17008" number="8" daytime="16:09" />
                <HEAT heatid="17009" number="9" daytime="16:10" />
                <HEAT heatid="17010" number="10" daytime="16:12" />
                <HEAT heatid="17011" number="11" daytime="16:13" />
                <HEAT heatid="17012" number="12" daytime="16:14" />
                <HEAT heatid="17013" number="13" daytime="16:15" />
                <HEAT heatid="17014" number="14" daytime="16:16" />
                <HEAT heatid="17015" number="15" daytime="16:18" />
                <HEAT heatid="17016" number="16" daytime="16:19" />
                <HEAT heatid="17017" number="17" daytime="16:20" />
                <HEAT heatid="17018" number="18" daytime="16:21" />
                <HEAT heatid="17019" number="19" daytime="16:22" />
                <HEAT heatid="17020" number="20" daytime="16:24" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="11" resultid="315" />
                    <RANKING place="13" resultid="396" />
                    <RANKING place="7" resultid="694" />
                    <RANKING place="4" resultid="865" />
                    <RANKING place="8" resultid="878" />
                    <RANKING place="6" resultid="896" />
                    <RANKING place="3" resultid="916" />
                    <RANKING place="15" resultid="1087" />
                    <RANKING place="9" resultid="1172" />
                    <RANKING place="2" resultid="1341" />
                    <RANKING place="5" resultid="1533" />
                    <RANKING place="12" resultid="1714" />
                    <RANKING place="14" resultid="1945" />
                    <RANKING place="10" resultid="1973" />
                    <RANKING place="1" resultid="2259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="1" resultid="18" />
                    <RANKING place="4" resultid="26" />
                    <RANKING place="10" resultid="39" />
                    <RANKING place="8" resultid="47" />
                    <RANKING place="6" resultid="51" />
                    <RANKING place="15" resultid="242" />
                    <RANKING place="11" resultid="565" />
                    <RANKING place="16" resultid="886" />
                    <RANKING place="14" resultid="1004" />
                    <RANKING place="2" resultid="1175" />
                    <RANKING place="9" resultid="1430" />
                    <RANKING place="7" resultid="1448" />
                    <RANKING place="5" resultid="1704" />
                    <RANKING place="12" resultid="1780" />
                    <RANKING place="13" resultid="2061" />
                    <RANKING place="3" resultid="2121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="6" resultid="210" />
                    <RANKING place="4" resultid="302" />
                    <RANKING place="2" resultid="345" />
                    <RANKING place="8" resultid="720" />
                    <RANKING place="9" resultid="1054" />
                    <RANKING place="7" resultid="1165" />
                    <RANKING place="1" resultid="1304" />
                    <RANKING place="12" resultid="1319" />
                    <RANKING place="10" resultid="1377" />
                    <RANKING place="11" resultid="1464" />
                    <RANKING place="3" resultid="1654" />
                    <RANKING place="5" resultid="1678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="8" resultid="80" />
                    <RANKING place="6" resultid="97" />
                    <RANKING place="7" resultid="118" />
                    <RANKING place="13" resultid="215" />
                    <RANKING place="2" resultid="350" />
                    <RANKING place="4" resultid="435" />
                    <RANKING place="11" resultid="892" />
                    <RANKING place="5" resultid="912" />
                    <RANKING place="12" resultid="1014" />
                    <RANKING place="3" resultid="1029" />
                    <RANKING place="10" resultid="1335" />
                    <RANKING place="1" resultid="1412" />
                    <RANKING place="9" resultid="1436" />
                    <RANKING place="15" resultid="1989" />
                    <RANKING place="14" resultid="2134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="104" />
                    <RANKING place="7" resultid="191" />
                    <RANKING place="3" resultid="249" />
                    <RANKING place="12" resultid="732" />
                    <RANKING place="8" resultid="984" />
                    <RANKING place="2" resultid="1187" />
                    <RANKING place="4" resultid="1309" />
                    <RANKING place="1" resultid="1480" />
                    <RANKING place="6" resultid="1570" />
                    <RANKING place="9" resultid="1888" />
                    <RANKING place="14" resultid="1967" />
                    <RANKING place="10" resultid="2009" />
                    <RANKING place="13" resultid="2227" />
                    <RANKING place="11" resultid="2234" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18" number="17" gender="M" round="TIM" order="17">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="18000" number="0" />
                <HEAT heatid="18001" number="1" daytime="16:28" />
                <HEAT heatid="18002" number="2" daytime="16:29" />
                <HEAT heatid="18003" number="3" daytime="16:31" />
                <HEAT heatid="18004" number="4" daytime="16:32" />
                <HEAT heatid="18005" number="5" daytime="16:34" />
                <HEAT heatid="18006" number="6" daytime="16:35" />
                <HEAT heatid="18007" number="7" daytime="16:36" />
                <HEAT heatid="18008" number="8" daytime="16:37" />
                <HEAT heatid="18009" number="9" daytime="16:38" />
                <HEAT heatid="18010" number="10" daytime="16:39" />
                <HEAT heatid="18011" number="11" daytime="16:41" />
                <HEAT heatid="18012" number="12" daytime="16:42" />
                <HEAT heatid="18013" number="13" daytime="16:43" />
                <HEAT heatid="18014" number="14" daytime="16:45" />
                <HEAT heatid="18015" number="15" daytime="16:46" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="2" resultid="376" />
                    <RANKING place="4" resultid="485" />
                    <RANKING place="5" resultid="1058" />
                    <RANKING place="3" resultid="1313" />
                    <RANKING place="1" resultid="1919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="10" resultid="22" />
                    <RANKING place="2" resultid="35" />
                    <RANKING place="8" resultid="221" />
                    <RANKING place="6" resultid="370" />
                    <RANKING place="7" resultid="588" />
                    <RANKING place="5" resultid="736" />
                    <RANKING place="9" resultid="754" />
                    <RANKING place="3" resultid="1700" />
                    <RANKING place="4" resultid="1755" />
                    <RANKING place="1" resultid="1985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="4" resultid="296" />
                    <RANKING place="3" resultid="670" />
                    <RANKING place="5" resultid="1000" />
                    <RANKING place="2" resultid="1795" />
                    <RANKING place="6" resultid="2162" />
                    <RANKING place="1" resultid="2254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="3" resultid="409" />
                    <RANKING place="1" resultid="962" />
                    <RANKING place="2" resultid="994" />
                    <RANKING place="5" resultid="1720" />
                    <RANKING place="4" resultid="2220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="76" />
                    <RANKING place="1" resultid="442" />
                    <RANKING place="2" resultid="1221" />
                    <RANKING place="8" resultid="1585" />
                    <RANKING place="6" resultid="1604" />
                    <RANKING place="7" resultid="1913" />
                    <RANKING place="3" resultid="2016" />
                    <RANKING place="4" resultid="2043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="266" />
                    <RANKING place="12" resultid="605" />
                    <RANKING place="11" resultid="726" />
                    <RANKING place="1" resultid="802" />
                    <RANKING place="4" resultid="1211" />
                    <RANKING place="6" resultid="1281" />
                    <RANKING place="2" resultid="1401" />
                    <RANKING place="13" resultid="1566" />
                    <RANKING place="7" resultid="1731" />
                    <RANKING place="5" resultid="1817" />
                    <RANKING place="9" resultid="1872" />
                    <RANKING place="10" resultid="1924" />
                    <RANKING place="8" resultid="1958" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="19" number="18" gender="F" round="TIM" order="18">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="19000" number="0" />
                <HEAT heatid="19001" number="1" daytime="16:50" />
                <HEAT heatid="19002" number="2" daytime="16:52" />
                <HEAT heatid="19003" number="3" daytime="16:55" />
                <HEAT heatid="19004" number="4" daytime="16:57" />
                <HEAT heatid="19005" number="5" daytime="17:00" />
                <HEAT heatid="19006" number="6" daytime="17:02" />
                <HEAT heatid="19007" number="7" daytime="17:04" />
                <HEAT heatid="19008" number="8" daytime="17:06" />
                <HEAT heatid="19009" number="9" daytime="17:08" />
                <HEAT heatid="19010" number="10" daytime="17:10" />
                <HEAT heatid="19011" number="11" daytime="17:12" />
                <HEAT heatid="19012" number="12" daytime="17:14" />
                <HEAT heatid="19013" number="13" daytime="17:16" />
                <HEAT heatid="19014" number="14" daytime="17:18" />
                <HEAT heatid="19015" number="15" daytime="17:20" />
                <HEAT heatid="19016" number="16" daytime="17:22" />
                <HEAT heatid="19017" number="17" daytime="17:23" />
                <HEAT heatid="19018" number="18" daytime="17:25" />
                <HEAT heatid="19019" number="19" daytime="17:27" />
                <HEAT heatid="19020" number="20" daytime="17:29" />
                <HEAT heatid="19021" number="21" daytime="17:30" />
                <HEAT heatid="19022" number="22" daytime="17:33" />
                <HEAT heatid="19023" number="23" daytime="17:34" />
                <HEAT heatid="19024" number="24" daytime="17:36" />
                <HEAT heatid="19025" number="25" daytime="17:38" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="8" resultid="316" />
                    <RANKING place="11" resultid="397" />
                    <RANKING place="5" resultid="456" />
                    <RANKING place="9" resultid="695" />
                    <RANKING place="7" resultid="866" />
                    <RANKING place="2" resultid="879" />
                    <RANKING place="1" resultid="897" />
                    <RANKING place="4" resultid="1342" />
                    <RANKING place="10" resultid="1534" />
                    <RANKING place="3" resultid="1555" />
                    <RANKING place="6" resultid="1715" />
                    <RANKING place="14" resultid="1900" />
                    <RANKING place="13" resultid="1946" />
                    <RANKING place="12" resultid="1974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="12" resultid="14" />
                    <RANKING place="5" resultid="19" />
                    <RANKING place="2" resultid="44" />
                    <RANKING place="18" resultid="243" />
                    <RANKING place="3" resultid="358" />
                    <RANKING place="4" resultid="502" />
                    <RANKING place="6" resultid="593" />
                    <RANKING place="9" resultid="701" />
                    <RANKING place="1" resultid="870" />
                    <RANKING place="19" resultid="887" />
                    <RANKING place="21" resultid="901" />
                    <RANKING place="14" resultid="1005" />
                    <RANKING place="7" resultid="1294" />
                    <RANKING place="10" resultid="1431" />
                    <RANKING place="13" resultid="1449" />
                    <RANKING place="11" resultid="1705" />
                    <RANKING place="16" resultid="1781" />
                    <RANKING place="15" resultid="1838" />
                    <RANKING place="20" resultid="2062" />
                    <RANKING place="17" resultid="2110" />
                    <RANKING place="8" resultid="2122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="9" resultid="303" />
                    <RANKING place="3" resultid="346" />
                    <RANKING place="5" resultid="721" />
                    <RANKING place="17" resultid="875" />
                    <RANKING place="10" resultid="1055" />
                    <RANKING place="4" resultid="1078" />
                    <RANKING place="1" resultid="1305" />
                    <RANKING place="12" resultid="1320" />
                    <RANKING place="14" resultid="1378" />
                    <RANKING place="13" resultid="1396" />
                    <RANKING place="18" resultid="1465" />
                    <RANKING place="6" resultid="1487" />
                    <RANKING place="15" resultid="1515" />
                    <RANKING place="2" resultid="1655" />
                    <RANKING place="11" resultid="1662" />
                    <RANKING place="8" resultid="1679" />
                    <RANKING place="7" resultid="1823" />
                    <RANKING place="16" resultid="2030" />
                    <RANKING place="19" resultid="2143" />
                    <RANKING place="20" resultid="2191" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="4" resultid="111" />
                    <RANKING place="7" resultid="119" />
                    <RANKING place="6" resultid="198" />
                    <RANKING place="9" resultid="204" />
                    <RANKING place="11" resultid="216" />
                    <RANKING place="1" resultid="255" />
                    <RANKING place="5" resultid="351" />
                    <RANKING place="8" resultid="436" />
                    <RANKING place="16" resultid="893" />
                    <RANKING place="14" resultid="1015" />
                    <RANKING place="17" resultid="1025" />
                    <RANKING place="10" resultid="1030" />
                    <RANKING place="2" resultid="1108" />
                    <RANKING place="13" resultid="1336" />
                    <RANKING place="12" resultid="1437" />
                    <RANKING place="3" resultid="1493" />
                    <RANKING place="15" resultid="1550" />
                    <RANKING place="18" resultid="2139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="12" resultid="105" />
                    <RANKING place="1" resultid="462" />
                    <RANKING place="9" resultid="522" />
                    <RANKING place="2" resultid="676" />
                    <RANKING place="5" resultid="733" />
                    <RANKING place="13" resultid="985" />
                    <RANKING place="10" resultid="1170" />
                    <RANKING place="3" resultid="1326" />
                    <RANKING place="7" resultid="1390" />
                    <RANKING place="4" resultid="1470" />
                    <RANKING place="14" resultid="1889" />
                    <RANKING place="16" resultid="1968" />
                    <RANKING place="11" resultid="2010" />
                    <RANKING place="6" resultid="2127" />
                    <RANKING place="15" resultid="2228" />
                    <RANKING place="8" resultid="2235" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="20" number="19" gender="M" round="TIM" order="19">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="20000" number="0" />
                <HEAT heatid="20001" number="1" daytime="17:42" />
                <HEAT heatid="20002" number="2" daytime="17:45" />
                <HEAT heatid="20003" number="3" daytime="17:47" />
                <HEAT heatid="20004" number="4" daytime="17:49" />
                <HEAT heatid="20005" number="5" daytime="17:52" />
                <HEAT heatid="20006" number="6" daytime="17:54" />
                <HEAT heatid="20007" number="7" daytime="17:56" />
                <HEAT heatid="20008" number="8" daytime="17:58" />
                <HEAT heatid="20009" number="9" daytime="18:00" />
                <HEAT heatid="20010" number="10" daytime="18:01" />
                <HEAT heatid="20011" number="11" daytime="18:03" />
                <HEAT heatid="20012" number="12" daytime="18:05" />
                <HEAT heatid="20013" number="13" daytime="18:07" />
                <HEAT heatid="20014" number="14" daytime="18:08" />
                <HEAT heatid="20015" number="15" daytime="18:10" />
                <HEAT heatid="20016" number="16" daytime="18:12" />
                <HEAT heatid="20017" number="17" daytime="18:13" />
                <HEAT heatid="20018" number="18" daytime="18:16" />
                <HEAT heatid="20019" number="19" daytime="18:17" />
                <HEAT heatid="20020" number="20" daytime="18:19" />
                <HEAT heatid="20021" number="21" daytime="18:21" />
                <HEAT heatid="20022" number="22" daytime="18:22" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2017">
                  <RANKINGS>
                    <RANKING place="4" resultid="473" />
                    <RANKING place="5" resultid="486" />
                    <RANKING place="2" resultid="528" />
                    <RANKING place="7" resultid="1059" />
                    <RANKING place="6" resultid="1314" />
                    <RANKING place="1" resultid="1630" />
                    <RANKING place="3" resultid="1920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2016">
                  <RANKINGS>
                    <RANKING place="2" resultid="5" />
                    <RANKING place="8" resultid="222" />
                    <RANKING place="1" resultid="327" />
                    <RANKING place="4" resultid="371" />
                    <RANKING place="6" resultid="589" />
                    <RANKING place="11" resultid="737" />
                    <RANKING place="13" resultid="755" />
                    <RANKING place="7" resultid="929" />
                    <RANKING place="3" resultid="1650" />
                    <RANKING place="5" resultid="1701" />
                    <RANKING place="10" resultid="1756" />
                    <RANKING place="12" resultid="1771" />
                    <RANKING place="9" resultid="1986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="10" resultid="232" />
                    <RANKING place="3" resultid="297" />
                    <RANKING place="5" resultid="422" />
                    <RANKING place="1" resultid="533" />
                    <RANKING place="7" resultid="671" />
                    <RANKING place="9" resultid="689" />
                    <RANKING place="6" resultid="1001" />
                    <RANKING place="8" resultid="1529" />
                    <RANKING place="2" resultid="1796" />
                    <RANKING place="11" resultid="2163" />
                    <RANKING place="4" resultid="2255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="10" resultid="290" />
                    <RANKING place="11" resultid="410" />
                    <RANKING place="1" resultid="548" />
                    <RANKING place="4" resultid="553" />
                    <RANKING place="9" resultid="939" />
                    <RANKING place="3" resultid="995" />
                    <RANKING place="2" resultid="1068" />
                    <RANKING place="7" resultid="1145" />
                    <RANKING place="6" resultid="1425" />
                    <RANKING place="12" resultid="1545" />
                    <RANKING place="15" resultid="1632" />
                    <RANKING place="5" resultid="1697" />
                    <RANKING place="14" resultid="1721" />
                    <RANKING place="8" resultid="1833" />
                    <RANKING place="13" resultid="1931" />
                    <RANKING place="17" resultid="2003" />
                    <RANKING place="16" resultid="2294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="7" resultid="10" />
                    <RANKING place="2" resultid="115" />
                    <RANKING place="5" resultid="186" />
                    <RANKING place="1" resultid="443" />
                    <RANKING place="8" resultid="512" />
                    <RANKING place="16" resultid="1083" />
                    <RANKING place="3" resultid="1222" />
                    <RANKING place="4" resultid="1442" />
                    <RANKING place="15" resultid="1586" />
                    <RANKING place="12" resultid="1605" />
                    <RANKING place="14" resultid="1914" />
                    <RANKING place="10" resultid="2017" />
                    <RANKING place="9" resultid="2044" />
                    <RANKING place="13" resultid="2051" />
                    <RANKING place="6" resultid="2068" />
                    <RANKING place="11" resultid="2157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="10" resultid="94" />
                    <RANKING place="4" resultid="267" />
                    <RANKING place="6" resultid="601" />
                    <RANKING place="9" resultid="727" />
                    <RANKING place="2" resultid="1212" />
                    <RANKING place="1" resultid="1282" />
                    <RANKING place="5" resultid="1402" />
                    <RANKING place="13" resultid="1567" />
                    <RANKING place="8" resultid="1732" />
                    <RANKING place="3" resultid="1818" />
                    <RANKING place="7" resultid="1873" />
                    <RANKING place="12" resultid="1925" />
                    <RANKING place="11" resultid="1959" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="21" number="20" gender="F" round="TIM" order="20">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="21001" number="1" daytime="18:27" />
                <HEAT heatid="21002" number="2" daytime="18:31" />
                <HEAT heatid="21003" number="3" daytime="18:35" />
                <HEAT heatid="21004" number="4" daytime="18:38" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="1" resultid="969" />
                    <RANKING place="3" resultid="1079" />
                    <RANKING place="2" resultid="1656" />
                    <RANKING place="4" resultid="1680" />
                    <RANKING place="5" resultid="1824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="112" />
                    <RANKING place="5" resultid="507" />
                    <RANKING place="3" resultid="1031" />
                    <RANKING place="4" resultid="1413" />
                    <RANKING place="2" resultid="1777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="192" />
                    <RANKING place="2" resultid="1232" />
                    <RANKING place="1" resultid="1481" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22" number="21" gender="M" round="TIM" order="21">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="22000" number="0" />
                <HEAT heatid="22002" number="2" daytime="18:49" />
                <HEAT heatid="22003" number="3" daytime="18:53" />
                <HEAT heatid="22004" number="4" daytime="18:57" />
                <HEAT heatid="22005" number="5" daytime="19:00" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="2" resultid="534" />
                    <RANKING place="1" resultid="1797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="5" resultid="291" />
                    <RANKING place="3" resultid="554" />
                    <RANKING place="4" resultid="560" />
                    <RANKING place="2" resultid="963" />
                    <RANKING place="1" resultid="1069" />
                    <RANKING place="6" resultid="1834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="444" />
                    <RANKING place="2" resultid="1443" />
                    <RANKING place="3" resultid="2069" />
                    <RANKING place="4" resultid="2158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="803" />
                    <RANKING place="3" resultid="1733" />
                    <RANKING place="2" resultid="2283" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23" number="22" gender="X" round="TIM" order="22">
              <SWIMSTYLE stroke="MEDLEY" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="23001" number="1" daytime="19:06" />
                <HEAT heatid="23002" number="2" daytime="19:09" />
                <HEAT heatid="23003" number="3" daytime="19:13" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="13" agemin="8" name="Jahrgänge 2012 bis 2017">
                  <RANKINGS>
                    <RANKING place="3" resultid="180" />
                    <RANKING place="2" resultid="280" />
                    <RANKING place="5" resultid="858" />
                    <RANKING place="7" resultid="859" />
                    <RANKING place="1" resultid="1288" />
                    <RANKING place="4" resultid="1850" />
                    <RANKING place="6" resultid="1856" />
                    <RANKING place="8" resultid="1862" />
                    <RANKING place="9" resultid="1866" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="3" date="2025-12-14" daytime="08:45" officialmeeting="08:15" warmupfrom="07:30">
          <EVENTS>
            <EVENT eventid="43" number="23" gender="F" round="PRE" order="23">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="43000" number="0" />
                <HEAT heatid="43001" number="1" daytime="08:45" />
                <HEAT heatid="43002" number="2" daytime="08:45" />
                <HEAT heatid="43003" number="3" daytime="08:46" />
                <HEAT heatid="43004" number="4" daytime="08:47" />
                <HEAT heatid="43005" number="5" daytime="08:48" />
                <HEAT heatid="43006" number="6" daytime="08:49" />
                <HEAT heatid="43007" number="7" daytime="08:50" />
                <HEAT heatid="43008" number="8" daytime="08:51" />
                <HEAT heatid="43009" number="9" daytime="08:52" />
                <HEAT heatid="43010" number="10" daytime="08:53" />
                <HEAT heatid="43011" number="11" daytime="08:54" />
                <HEAT heatid="43012" number="12" daytime="08:55" />
                <HEAT heatid="43013" number="13" daytime="08:55" />
                <HEAT heatid="43014" number="14" daytime="08:56" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="9" resultid="57" />
                    <RANKING place="10" resultid="64" />
                    <RANKING place="3" resultid="223" />
                    <RANKING place="2" resultid="359" />
                    <RANKING place="6" resultid="474" />
                    <RANKING place="1" resultid="1352" />
                    <RANKING place="7" resultid="1663" />
                    <RANKING place="4" resultid="1736" />
                    <RANKING place="8" resultid="2031" />
                    <RANKING place="5" resultid="2094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="5" resultid="123" />
                    <RANKING place="6" resultid="167" />
                    <RANKING place="1" resultid="328" />
                    <RANKING place="8" resultid="637" />
                    <RANKING place="2" resultid="769" />
                    <RANKING place="9" resultid="1166" />
                    <RANKING place="10" resultid="1176" />
                    <RANKING place="3" resultid="1243" />
                    <RANKING place="7" resultid="1559" />
                    <RANKING place="4" resultid="2087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="20" resultid="141" />
                    <RANKING place="17" resultid="158" />
                    <RANKING place="5" resultid="377" />
                    <RANKING place="12" resultid="411" />
                    <RANKING place="24" resultid="611" />
                    <RANKING place="9" resultid="617" />
                    <RANKING place="12" resultid="621" />
                    <RANKING place="10" resultid="644" />
                    <RANKING place="7" resultid="678" />
                    <RANKING place="1" resultid="702" />
                    <RANKING place="11" resultid="831" />
                    <RANKING place="8" resultid="1109" />
                    <RANKING place="2" resultid="1122" />
                    <RANKING place="6" resultid="1193" />
                    <RANKING place="14" resultid="1203" />
                    <RANKING place="15" resultid="1223" />
                    <RANKING place="19" resultid="1233" />
                    <RANKING place="21" resultid="1253" />
                    <RANKING place="3" resultid="1263" />
                    <RANKING place="4" resultid="1379" />
                    <RANKING place="16" resultid="1450" />
                    <RANKING place="23" resultid="1597" />
                    <RANKING place="18" resultid="1947" />
                    <RANKING place="22" resultid="2053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="4" resultid="154" />
                    <RANKING place="1" resultid="818" />
                    <RANKING place="2" resultid="1041" />
                    <RANKING place="5" resultid="1571" />
                    <RANKING place="3" resultid="2176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="274" />
                    <RANKING place="3" resultid="1587" />
                    <RANKING place="1" resultid="2170" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="44" number="24" gender="M" round="PRE" order="24">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="44000" number="0" />
                <HEAT heatid="44001" number="1" daytime="08:59" />
                <HEAT heatid="44002" number="2" daytime="09:00" />
                <HEAT heatid="44003" number="3" daytime="09:01" />
                <HEAT heatid="44004" number="4" daytime="09:02" />
                <HEAT heatid="44005" number="5" daytime="09:03" />
                <HEAT heatid="44006" number="6" daytime="09:04" />
                <HEAT heatid="44007" number="7" daytime="09:05" />
                <HEAT heatid="44008" number="8" daytime="09:05" />
                <HEAT heatid="44009" number="9" daytime="09:06" />
                <HEAT heatid="44010" number="10" daytime="09:07" />
                <HEAT heatid="44011" number="11" daytime="09:08" />
                <HEAT heatid="44012" number="12" daytime="09:09" />
                <HEAT heatid="44013" number="13" daytime="09:09" />
                <HEAT heatid="44014" number="14" daytime="09:10" />
                <HEAT heatid="44015" number="15" daytime="09:11" />
                <HEAT heatid="44016" number="16" daytime="09:12" />
                <HEAT heatid="44017" number="17" daytime="09:13" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="9" resultid="120" />
                    <RANKING place="11" resultid="256" />
                    <RANKING place="7" resultid="626" />
                    <RANKING place="3" resultid="659" />
                    <RANKING place="1" resultid="1213" />
                    <RANKING place="8" resultid="1273" />
                    <RANKING place="5" resultid="1500" />
                    <RANKING place="12" resultid="1611" />
                    <RANKING place="6" resultid="1669" />
                    <RANKING place="10" resultid="1876" />
                    <RANKING place="2" resultid="1890" />
                    <RANKING place="4" resultid="2284" />
                    <RANKING place="13" resultid="2295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="11" resultid="61" />
                    <RANKING place="12" resultid="132" />
                    <RANKING place="5" resultid="145" />
                    <RANKING place="14" resultid="268" />
                    <RANKING place="7" resultid="493" />
                    <RANKING place="20" resultid="513" />
                    <RANKING place="24" resultid="631" />
                    <RANKING place="8" resultid="650" />
                    <RANKING place="19" resultid="773" />
                    <RANKING place="13" resultid="784" />
                    <RANKING place="10" resultid="810" />
                    <RANKING place="23" resultid="814" />
                    <RANKING place="6" resultid="1032" />
                    <RANKING place="22" resultid="1060" />
                    <RANKING place="1" resultid="1113" />
                    <RANKING place="9" resultid="1127" />
                    <RANKING place="2" resultid="1136" />
                    <RANKING place="26" resultid="1238" />
                    <RANKING place="18" resultid="1248" />
                    <RANKING place="21" resultid="1346" />
                    <RANKING place="29" resultid="1606" />
                    <RANKING place="4" resultid="1687" />
                    <RANKING place="3" resultid="1722" />
                    <RANKING place="15" resultid="1742" />
                    <RANKING place="28" resultid="1901" />
                    <RANKING place="25" resultid="1934" />
                    <RANKING place="16" resultid="2100" />
                    <RANKING place="27" resultid="2205" />
                    <RANKING place="17" resultid="2242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="1" resultid="385" />
                    <RANKING place="4" resultid="423" />
                    <RANKING place="2" resultid="445" />
                    <RANKING place="5" resultid="777" />
                    <RANKING place="9" resultid="796" />
                    <RANKING place="6" resultid="948" />
                    <RANKING place="3" resultid="1094" />
                    <RANKING place="8" resultid="1258" />
                    <RANKING place="7" resultid="1327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="463" />
                    <RANKING place="6" resultid="804" />
                    <RANKING place="5" resultid="843" />
                    <RANKING place="3" resultid="1160" />
                    <RANKING place="7" resultid="1343" />
                    <RANKING place="10" resultid="1414" />
                    <RANKING place="4" resultid="1456" />
                    <RANKING place="9" resultid="1521" />
                    <RANKING place="8" resultid="1592" />
                    <RANKING place="1" resultid="2148" />
                    <RANKING place="11" resultid="2266" />
                    <RANKING place="12" resultid="2268" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="27" number="25" gender="F" round="PRE" order="25">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="27000" number="0" />
                <HEAT heatid="27001" number="1" daytime="09:15" />
                <HEAT heatid="27002" number="2" daytime="09:17" />
                <HEAT heatid="27003" number="3" daytime="09:18" />
                <HEAT heatid="27004" number="4" daytime="09:19" />
                <HEAT heatid="27005" number="5" daytime="09:20" />
                <HEAT heatid="27006" number="6" daytime="09:21" />
                <HEAT heatid="27007" number="7" daytime="09:22" />
                <HEAT heatid="27008" number="8" daytime="09:23" />
                <HEAT heatid="27009" number="9" daytime="09:24" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="58" />
                    <RANKING place="9" resultid="65" />
                    <RANKING place="8" resultid="224" />
                    <RANKING place="6" resultid="475" />
                    <RANKING place="1" resultid="1353" />
                    <RANKING place="4" resultid="1664" />
                    <RANKING place="5" resultid="2032" />
                    <RANKING place="7" resultid="2095" />
                    <RANKING place="3" resultid="2274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="7" resultid="99" />
                    <RANKING place="5" resultid="168" />
                    <RANKING place="3" resultid="329" />
                    <RANKING place="6" resultid="638" />
                    <RANKING place="9" resultid="1167" />
                    <RANKING place="1" resultid="1244" />
                    <RANKING place="4" resultid="1560" />
                    <RANKING place="2" resultid="1975" />
                    <RANKING place="8" resultid="2182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="13" resultid="159" />
                    <RANKING place="8" resultid="334" />
                    <RANKING place="9" resultid="622" />
                    <RANKING place="10" resultid="645" />
                    <RANKING place="2" resultid="679" />
                    <RANKING place="6" resultid="832" />
                    <RANKING place="4" resultid="1099" />
                    <RANKING place="1" resultid="1123" />
                    <RANKING place="5" resultid="1194" />
                    <RANKING place="11" resultid="1254" />
                    <RANKING place="7" resultid="1264" />
                    <RANKING place="3" resultid="1380" />
                    <RANKING place="12" resultid="1598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="2" resultid="788" />
                    <RANKING place="3" resultid="1572" />
                    <RANKING place="1" resultid="1706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="847" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="28" number="26" gender="M" round="PRE" order="26">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="28000" number="0" />
                <HEAT heatid="28001" number="1" daytime="09:27" />
                <HEAT heatid="28002" number="2" daytime="09:28" />
                <HEAT heatid="28003" number="3" daytime="09:29" />
                <HEAT heatid="28004" number="4" daytime="09:30" />
                <HEAT heatid="28005" number="5" daytime="09:31" />
                <HEAT heatid="28006" number="6" daytime="09:32" />
                <HEAT heatid="28007" number="7" daytime="09:33" />
                <HEAT heatid="28008" number="8" daytime="09:34" />
                <HEAT heatid="28009" number="9" daytime="09:35" />
                <HEAT heatid="28010" number="10" daytime="09:36" />
                <HEAT heatid="28011" number="11" daytime="09:37" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="9" resultid="257" />
                    <RANKING place="4" resultid="660" />
                    <RANKING place="2" resultid="766" />
                    <RANKING place="1" resultid="1188" />
                    <RANKING place="8" resultid="1198" />
                    <RANKING place="3" resultid="1214" />
                    <RANKING place="5" resultid="1274" />
                    <RANKING place="7" resultid="1501" />
                    <RANKING place="10" resultid="1612" />
                    <RANKING place="6" resultid="1877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="12" resultid="82" />
                    <RANKING place="5" resultid="146" />
                    <RANKING place="9" resultid="269" />
                    <RANKING place="7" resultid="535" />
                    <RANKING place="13" resultid="632" />
                    <RANKING place="6" resultid="651" />
                    <RANKING place="8" resultid="940" />
                    <RANKING place="4" resultid="944" />
                    <RANKING place="3" resultid="970" />
                    <RANKING place="2" resultid="1114" />
                    <RANKING place="1" resultid="1118" />
                    <RANKING place="11" resultid="1347" />
                    <RANKING place="16" resultid="1607" />
                    <RANKING place="15" resultid="1902" />
                    <RANKING place="10" resultid="1935" />
                    <RANKING place="14" resultid="2206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="5" resultid="85" />
                    <RANKING place="1" resultid="424" />
                    <RANKING place="2" resultid="778" />
                    <RANKING place="3" resultid="837" />
                    <RANKING place="4" resultid="1259" />
                    <RANKING place="6" resultid="2019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="655" />
                    <RANKING place="8" resultid="682" />
                    <RANKING place="1" resultid="807" />
                    <RANKING place="3" resultid="844" />
                    <RANKING place="7" resultid="1344" />
                    <RANKING place="2" resultid="1360" />
                    <RANKING place="5" resultid="1415" />
                    <RANKING place="6" resultid="2267" />
                    <RANKING place="9" resultid="2269" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="29" number="27" gender="F" round="TIM" order="27">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="29000" number="0" />
                <HEAT heatid="29001" number="1" daytime="09:40" />
                <HEAT heatid="29002" number="2" daytime="09:42" />
                <HEAT heatid="29003" number="3" daytime="09:44" />
                <HEAT heatid="29004" number="4" daytime="09:45" />
                <HEAT heatid="29005" number="5" daytime="09:47" />
                <HEAT heatid="29006" number="6" daytime="09:49" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="360" />
                    <RANKING place="3" resultid="1354" />
                    <RANKING place="4" resultid="1737" />
                    <RANKING place="1" resultid="1798" />
                    <RANKING place="5" resultid="2275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="487" />
                    <RANKING place="1" resultid="1976" />
                    <RANKING place="2" resultid="2088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="6" resultid="335" />
                    <RANKING place="1" resultid="378" />
                    <RANKING place="5" resultid="412" />
                    <RANKING place="2" resultid="618" />
                    <RANKING place="4" resultid="1204" />
                    <RANKING place="8" resultid="1234" />
                    <RANKING place="3" resultid="1839" />
                    <RANKING place="7" resultid="2054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="1" resultid="1131" />
                    <RANKING place="2" resultid="1356" />
                    <RANKING place="3" resultid="2177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="1506" />
                    <RANKING place="1" resultid="2171" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="30" number="28" gender="M" round="TIM" order="28">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="30000" number="0" />
                <HEAT heatid="30001" number="1" daytime="09:53" />
                <HEAT heatid="30002" number="2" daytime="09:54" />
                <HEAT heatid="30003" number="3" daytime="09:56" />
                <HEAT heatid="30004" number="4" daytime="09:58" />
                <HEAT heatid="30005" number="5" daytime="09:59" />
                <HEAT heatid="30006" number="6" daytime="10:00" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="1891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="10" resultid="106" />
                    <RANKING place="7" resultid="133" />
                    <RANKING place="8" resultid="514" />
                    <RANKING place="4" resultid="811" />
                    <RANKING place="5" resultid="1006" />
                    <RANKING place="2" resultid="1033" />
                    <RANKING place="11" resultid="1249" />
                    <RANKING place="1" resultid="1688" />
                    <RANKING place="3" resultid="1723" />
                    <RANKING place="6" resultid="1743" />
                    <RANKING place="9" resultid="2243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="386" />
                    <RANKING place="2" resultid="446" />
                    <RANKING place="4" resultid="838" />
                    <RANKING place="1" resultid="1095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="464" />
                    <RANKING place="4" resultid="793" />
                    <RANKING place="3" resultid="1156" />
                    <RANKING place="2" resultid="1361" />
                    <RANKING place="5" resultid="1416" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="47" number="29" gender="F" round="TIM" order="29">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="47000" number="0" />
                <HEAT heatid="47001" number="1" daytime="10:04" />
                <HEAT heatid="47002" number="2" daytime="10:06" />
                <HEAT heatid="47003" number="3" daytime="10:08" />
                <HEAT heatid="47004" number="4" daytime="10:10" />
                <HEAT heatid="47005" number="5" daytime="10:12" />
                <HEAT heatid="47006" number="6" daytime="10:14" />
                <HEAT heatid="47007" number="7" daytime="10:15" />
                <HEAT heatid="47008" number="8" daytime="10:17" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="476" />
                    <RANKING place="5" resultid="540" />
                    <RANKING place="2" resultid="1738" />
                    <RANKING place="1" resultid="1799" />
                    <RANKING place="4" resultid="2033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="124" />
                    <RANKING place="1" resultid="330" />
                    <RANKING place="3" resultid="488" />
                    <RANKING place="5" resultid="1177" />
                    <RANKING place="4" resultid="2183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="10" resultid="142" />
                    <RANKING place="3" resultid="379" />
                    <RANKING place="6" resultid="646" />
                    <RANKING place="4" resultid="780" />
                    <RANKING place="1" resultid="1110" />
                    <RANKING place="9" resultid="1224" />
                    <RANKING place="11" resultid="1255" />
                    <RANKING place="2" resultid="1381" />
                    <RANKING place="7" resultid="1451" />
                    <RANKING place="5" resultid="1840" />
                    <RANKING place="8" resultid="1948" />
                    <RANKING place="12" resultid="2055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="1" resultid="1042" />
                    <RANKING place="2" resultid="1357" />
                    <RANKING place="3" resultid="2178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="1507" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="48" number="30" gender="M" round="TIM" order="30">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="48000" number="0" />
                <HEAT heatid="48001" number="1" daytime="10:21" />
                <HEAT heatid="48002" number="2" daytime="10:23" />
                <HEAT heatid="48003" number="3" daytime="10:24" />
                <HEAT heatid="48004" number="4" daytime="10:26" />
                <HEAT heatid="48005" number="5" daytime="10:27" />
                <HEAT heatid="48006" number="6" daytime="10:29" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="138" />
                    <RANKING place="5" resultid="258" />
                    <RANKING place="4" resultid="1275" />
                    <RANKING place="3" resultid="1892" />
                    <RANKING place="1" resultid="2285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="3" resultid="515" />
                    <RANKING place="4" resultid="774" />
                    <RANKING place="1" resultid="1007" />
                    <RANKING place="2" resultid="1128" />
                    <RANKING place="6" resultid="1239" />
                    <RANKING place="7" resultid="1903" />
                    <RANKING place="5" resultid="2244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="2" resultid="425" />
                    <RANKING place="4" resultid="797" />
                    <RANKING place="1" resultid="949" />
                    <RANKING place="3" resultid="1328" />
                    <RANKING place="5" resultid="2020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="1522" />
                    <RANKING place="1" resultid="1593" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="33" number="31" gender="F" round="TIM" order="31">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="33000" number="0" />
                <HEAT heatid="33001" number="1" daytime="10:32" />
                <HEAT heatid="33002" number="2" daytime="10:35" />
                <HEAT heatid="33003" number="3" daytime="10:37" />
                <HEAT heatid="33004" number="4" daytime="10:38" />
                <HEAT heatid="33005" number="5" daytime="10:40" />
                <HEAT heatid="33006" number="6" daytime="10:42" />
                <HEAT heatid="33007" number="7" daytime="10:44" />
                <HEAT heatid="33008" number="8" daytime="10:45" />
                <HEAT heatid="33009" number="9" daytime="10:47" />
                <HEAT heatid="33010" number="10" daytime="10:49" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="361" />
                    <RANKING place="6" resultid="541" />
                    <RANKING place="1" resultid="1355" />
                    <RANKING place="3" resultid="1800" />
                    <RANKING place="5" resultid="2034" />
                    <RANKING place="4" resultid="2096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="169" />
                    <RANKING place="5" resultid="489" />
                    <RANKING place="7" resultid="639" />
                    <RANKING place="1" resultid="770" />
                    <RANKING place="2" resultid="1245" />
                    <RANKING place="8" resultid="1561" />
                    <RANKING place="3" resultid="1977" />
                    <RANKING place="4" resultid="2089" />
                    <RANKING place="9" resultid="2184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="8" resultid="336" />
                    <RANKING place="5" resultid="380" />
                    <RANKING place="9" resultid="413" />
                    <RANKING place="12" resultid="613" />
                    <RANKING place="2" resultid="1100" />
                    <RANKING place="1" resultid="1124" />
                    <RANKING place="3" resultid="1195" />
                    <RANKING place="10" resultid="1235" />
                    <RANKING place="6" resultid="1265" />
                    <RANKING place="4" resultid="1382" />
                    <RANKING place="11" resultid="1599" />
                    <RANKING place="6" resultid="1841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="155" />
                    <RANKING place="2" resultid="789" />
                    <RANKING place="4" resultid="1573" />
                    <RANKING place="1" resultid="1707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="126" />
                    <RANKING place="2" resultid="275" />
                    <RANKING place="3" resultid="1588" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="34" number="32" gender="M" round="TIM" order="32">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="34000" number="0" />
                <HEAT heatid="34001" number="1" daytime="10:52" />
                <HEAT heatid="34002" number="2" daytime="10:54" />
                <HEAT heatid="34003" number="3" daytime="10:56" />
                <HEAT heatid="34004" number="4" daytime="10:58" />
                <HEAT heatid="34005" number="5" daytime="11:00" />
                <HEAT heatid="34006" number="6" daytime="11:01" />
                <HEAT heatid="34007" number="7" daytime="11:03" />
                <HEAT heatid="34008" number="8" daytime="11:04" />
                <HEAT heatid="34009" number="9" daytime="11:06" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="9" resultid="121" />
                    <RANKING place="6" resultid="628" />
                    <RANKING place="3" resultid="661" />
                    <RANKING place="1" resultid="1189" />
                    <RANKING place="7" resultid="1199" />
                    <RANKING place="2" resultid="1215" />
                    <RANKING place="5" resultid="1502" />
                    <RANKING place="4" resultid="1670" />
                    <RANKING place="8" resultid="1878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="10" resultid="83" />
                    <RANKING place="9" resultid="107" />
                    <RANKING place="2" resultid="147" />
                    <RANKING place="13" resultid="174" />
                    <RANKING place="5" resultid="270" />
                    <RANKING place="4" resultid="494" />
                    <RANKING place="3" resultid="536" />
                    <RANKING place="12" resultid="633" />
                    <RANKING place="8" resultid="1061" />
                    <RANKING place="1" resultid="1115" />
                    <RANKING place="6" resultid="1250" />
                    <RANKING place="7" resultid="1744" />
                    <RANKING place="11" resultid="1936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="86" />
                    <RANKING place="1" resultid="387" />
                    <RANKING place="2" resultid="1329" />
                    <RANKING place="4" resultid="2021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="805" />
                    <RANKING place="5" resultid="1157" />
                    <RANKING place="1" resultid="1362" />
                    <RANKING place="2" resultid="1457" />
                    <RANKING place="3" resultid="1471" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="51" number="33" gender="F" round="TIM" order="33">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="51000" number="0" />
                <HEAT heatid="51001" number="1" daytime="11:09" />
                <HEAT heatid="51002" number="2" daytime="11:13" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="781" />
                    <RANKING place="1" resultid="819" />
                    <RANKING place="4" resultid="1452" />
                    <RANKING place="6" resultid="1665" />
                    <RANKING place="5" resultid="1949" />
                    <RANKING place="7" resultid="2128" />
                    <RANKING place="2" resultid="2172" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="52" number="34" gender="M" round="TIM" order="34">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="52000" number="0" />
                <HEAT heatid="52001" number="1" daytime="11:16" />
                <HEAT heatid="52002" number="2" daytime="11:19" />
                <HEAT heatid="52003" number="3" daytime="11:22" />
                <HEAT heatid="52004" number="4" daytime="11:25" />
                <HEAT heatid="52005" number="5" daytime="11:28" />
                <HEAT heatid="52006" number="6" daytime="11:31" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="8" resultid="134" />
                    <RANKING place="2" resultid="388" />
                    <RANKING place="9" resultid="495" />
                    <RANKING place="16" resultid="634" />
                    <RANKING place="15" resultid="662" />
                    <RANKING place="10" resultid="785" />
                    <RANKING place="6" resultid="794" />
                    <RANKING place="14" resultid="815" />
                    <RANKING place="4" resultid="1034" />
                    <RANKING place="3" resultid="1137" />
                    <RANKING place="12" resultid="1348" />
                    <RANKING place="1" resultid="1363" />
                    <RANKING place="13" resultid="1671" />
                    <RANKING place="7" resultid="1689" />
                    <RANKING place="5" resultid="1724" />
                    <RANKING place="18" resultid="1874" />
                    <RANKING place="21" resultid="1932" />
                    <RANKING place="20" resultid="2052" />
                    <RANKING place="17" resultid="2070" />
                    <RANKING place="19" resultid="2208" />
                    <RANKING place="11" resultid="2245" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="37" number="35" gender="F" round="TIM" order="35">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="37000" number="0" />
                <HEAT heatid="37001" number="1" daytime="11:33" />
                <HEAT heatid="37002" number="2" daytime="11:37" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="59" />
                    <RANKING place="8" resultid="81" />
                    <RANKING place="7" resultid="98" />
                    <RANKING place="4" resultid="337" />
                    <RANKING place="1" resultid="523" />
                    <RANKING place="3" resultid="1132" />
                    <RANKING place="2" resultid="1708" />
                    <RANKING place="5" resultid="2276" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="38" number="36" gender="M" round="TIM" order="36">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="38000" number="0" />
                <HEAT heatid="38001" number="1" daytime="11:42" />
                <HEAT heatid="38002" number="2" daytime="11:47" />
                <HEAT heatid="38003" number="3" daytime="11:51" />
                <HEAT heatid="38004" number="4" daytime="11:55" />
                <HEAT heatid="38005" number="5" daytime="11:58" />
                <HEAT heatid="38006" number="6" daytime="12:01" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="19" resultid="77" />
                    <RANKING place="5" resultid="426" />
                    <RANKING place="9" resultid="537" />
                    <RANKING place="8" resultid="652" />
                    <RANKING place="12" resultid="767" />
                    <RANKING place="6" resultid="839" />
                    <RANKING place="7" resultid="941" />
                    <RANKING place="3" resultid="945" />
                    <RANKING place="2" resultid="971" />
                    <RANKING place="1" resultid="1119" />
                    <RANKING place="10" resultid="1190" />
                    <RANKING place="11" resultid="1349" />
                    <RANKING place="4" resultid="1472" />
                    <RANKING place="14" resultid="1503" />
                    <RANKING place="15" resultid="1734" />
                    <RANKING place="13" resultid="1879" />
                    <RANKING place="20" resultid="1904" />
                    <RANKING place="21" resultid="1915" />
                    <RANKING place="16" resultid="2018" />
                    <RANKING place="18" resultid="2045" />
                    <RANKING place="22" resultid="2221" />
                    <RANKING place="17" resultid="2256" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="39" number="37" gender="F" round="TIM" order="37">
              <SWIMSTYLE stroke="FREE" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="39001" number="1" daytime="12:06" />
                <HEAT heatid="39002" number="2" daytime="12:09" />
                <HEAT heatid="39003" number="3" daytime="12:11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Jahrgänge 2015 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="281" />
                    <RANKING place="5" resultid="608" />
                    <RANKING place="4" resultid="764" />
                    <RANKING place="1" resultid="860" />
                    <RANKING place="2" resultid="1178" />
                    <RANKING place="6" resultid="1285" />
                    <RANKING place="7" resultid="1847" />
                    <RANKING place="8" resultid="1853" />
                    <RANKING place="9" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="40" number="38" gender="M" round="TIM" order="38">
              <SWIMSTYLE stroke="FREE" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="40001" number="1" daytime="12:16" />
                <HEAT heatid="40002" number="2" daytime="12:18" />
                <HEAT heatid="40003" number="3" daytime="12:21" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Jahrgänge 2015 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="282" />
                    <RANKING place="4" resultid="606" />
                    <RANKING place="3" resultid="762" />
                    <RANKING place="6" resultid="862" />
                    <RANKING place="7" resultid="1180" />
                    <RANKING place="1" resultid="1283" />
                    <RANKING place="4" resultid="1845" />
                    <RANKING place="8" resultid="1851" />
                    <RANKING place="9" resultid="1857" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="4" date="2025-12-14" daytime="00:30">
          <EVENTS>
            <EVENT eventid="41" number="39" gender="F" round="PRE" order="39">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="41000" number="0" />
                <HEAT heatid="41001" number="1" daytime="12:55" />
                <HEAT heatid="41002" number="2" daytime="12:56" />
                <HEAT heatid="41003" number="3" daytime="12:57" />
                <HEAT heatid="41004" number="4" daytime="12:58" />
                <HEAT heatid="41005" number="5" daytime="12:59" />
                <HEAT heatid="41006" number="6" daytime="13:00" />
                <HEAT heatid="41007" number="7" daytime="13:01" />
                <HEAT heatid="41008" number="8" daytime="13:02" />
                <HEAT heatid="41009" number="9" daytime="13:03" />
                <HEAT heatid="41010" number="10" daytime="13:04" />
                <HEAT heatid="41011" number="11" daytime="13:04" />
                <HEAT heatid="41012" number="12" daytime="13:05" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="225" />
                    <RANKING place="1" resultid="362" />
                    <RANKING place="6" resultid="477" />
                    <RANKING place="5" resultid="1666" />
                    <RANKING place="2" resultid="1739" />
                    <RANKING place="7" resultid="2035" />
                    <RANKING place="4" resultid="2097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="490" />
                    <RANKING place="5" resultid="640" />
                    <RANKING place="1" resultid="771" />
                    <RANKING place="7" resultid="1562" />
                    <RANKING place="2" resultid="1978" />
                    <RANKING place="3" resultid="2090" />
                    <RANKING place="6" resultid="2185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="16" resultid="338" />
                    <RANKING place="4" resultid="381" />
                    <RANKING place="11" resultid="414" />
                    <RANKING place="21" resultid="614" />
                    <RANKING place="7" resultid="619" />
                    <RANKING place="18" resultid="623" />
                    <RANKING place="12" resultid="647" />
                    <RANKING place="9" resultid="680" />
                    <RANKING place="1" resultid="703" />
                    <RANKING place="5" resultid="1101" />
                    <RANKING place="2" resultid="1125" />
                    <RANKING place="6" resultid="1196" />
                    <RANKING place="14" resultid="1206" />
                    <RANKING place="15" resultid="1225" />
                    <RANKING place="20" resultid="1236" />
                    <RANKING place="17" resultid="1256" />
                    <RANKING place="8" resultid="1266" />
                    <RANKING place="3" resultid="1383" />
                    <RANKING place="13" resultid="1453" />
                    <RANKING place="10" resultid="1842" />
                    <RANKING place="19" resultid="2056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="4" resultid="156" />
                    <RANKING place="3" resultid="790" />
                    <RANKING place="1" resultid="1133" />
                    <RANKING place="5" resultid="1574" />
                    <RANKING place="2" resultid="2179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="127" />
                    <RANKING place="4" resultid="276" />
                    <RANKING place="3" resultid="1589" />
                    <RANKING place="1" resultid="2173" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="42" number="40" gender="M" round="PRE" order="40">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="42000" number="0" />
                <HEAT heatid="42001" number="1" daytime="13:08" />
                <HEAT heatid="42002" number="2" daytime="13:09" />
                <HEAT heatid="42003" number="3" daytime="13:10" />
                <HEAT heatid="42004" number="4" daytime="13:11" />
                <HEAT heatid="42005" number="5" daytime="13:12" />
                <HEAT heatid="42006" number="6" daytime="13:13" />
                <HEAT heatid="42007" number="7" daytime="13:14" />
                <HEAT heatid="42008" number="8" daytime="13:15" />
                <HEAT heatid="42009" number="9" daytime="13:16" />
                <HEAT heatid="42010" number="10" daytime="13:16" />
                <HEAT heatid="42011" number="11" daytime="13:17" />
                <HEAT heatid="42012" number="12" daytime="13:18" />
                <HEAT heatid="42013" number="13" daytime="13:19" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="5" resultid="629" />
                    <RANKING place="3" resultid="663" />
                    <RANKING place="6" resultid="1200" />
                    <RANKING place="4" resultid="1216" />
                    <RANKING place="7" resultid="1276" />
                    <RANKING place="9" resultid="1613" />
                    <RANKING place="2" resultid="1672" />
                    <RANKING place="8" resultid="1880" />
                    <RANKING place="1" resultid="1893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="11" resultid="62" />
                    <RANKING place="8" resultid="148" />
                    <RANKING place="14" resultid="271" />
                    <RANKING place="9" resultid="496" />
                    <RANKING place="6" resultid="516" />
                    <RANKING place="18" resultid="635" />
                    <RANKING place="10" resultid="653" />
                    <RANKING place="13" resultid="786" />
                    <RANKING place="6" resultid="812" />
                    <RANKING place="15" resultid="816" />
                    <RANKING place="5" resultid="1035" />
                    <RANKING place="17" resultid="1062" />
                    <RANKING place="1" resultid="1116" />
                    <RANKING place="3" resultid="1138" />
                    <RANKING place="20" resultid="1240" />
                    <RANKING place="21" resultid="1608" />
                    <RANKING place="2" resultid="1690" />
                    <RANKING place="4" resultid="1725" />
                    <RANKING place="12" resultid="1745" />
                    <RANKING place="19" resultid="1937" />
                    <RANKING place="16" resultid="2246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="389" />
                    <RANKING place="5" resultid="427" />
                    <RANKING place="2" resultid="447" />
                    <RANKING place="4" resultid="840" />
                    <RANKING place="1" resultid="1096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="465" />
                    <RANKING place="12" resultid="656" />
                    <RANKING place="9" resultid="795" />
                    <RANKING place="4" resultid="845" />
                    <RANKING place="7" resultid="1158" />
                    <RANKING place="5" resultid="1161" />
                    <RANKING place="10" resultid="1345" />
                    <RANKING place="6" resultid="1364" />
                    <RANKING place="11" resultid="1417" />
                    <RANKING place="2" resultid="1458" />
                    <RANKING place="8" resultid="1594" />
                    <RANKING place="1" resultid="2150" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="25" number="41" gender="F" round="PRE" order="41">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="25000" number="0" />
                <HEAT heatid="25001" number="1" daytime="13:22" />
                <HEAT heatid="25002" number="2" daytime="13:23" />
                <HEAT heatid="25003" number="3" daytime="13:24" />
                <HEAT heatid="25004" number="4" daytime="13:25" />
                <HEAT heatid="25005" number="5" daytime="13:26" />
                <HEAT heatid="25006" number="6" daytime="13:27" />
                <HEAT heatid="25007" number="7" daytime="13:28" />
                <HEAT heatid="25008" number="8" daytime="13:29" />
                <HEAT heatid="25009" number="9" daytime="13:30" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="5" resultid="66" />
                    <RANKING place="3" resultid="226" />
                    <RANKING place="1" resultid="363" />
                    <RANKING place="4" resultid="478" />
                    <RANKING place="7" resultid="542" />
                    <RANKING place="2" resultid="1801" />
                    <RANKING place="6" resultid="2036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="331" />
                    <RANKING place="4" resultid="491" />
                    <RANKING place="1" resultid="1246" />
                    <RANKING place="3" resultid="2091" />
                    <RANKING place="5" resultid="2186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="13" resultid="143" />
                    <RANKING place="11" resultid="160" />
                    <RANKING place="4" resultid="382" />
                    <RANKING place="10" resultid="415" />
                    <RANKING place="12" resultid="615" />
                    <RANKING place="6" resultid="648" />
                    <RANKING place="5" resultid="681" />
                    <RANKING place="1" resultid="704" />
                    <RANKING place="7" resultid="782" />
                    <RANKING place="3" resultid="1111" />
                    <RANKING place="9" resultid="1226" />
                    <RANKING place="2" resultid="1384" />
                    <RANKING place="8" resultid="1950" />
                    <RANKING place="14" resultid="2057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="1" resultid="1043" />
                    <RANKING place="2" resultid="2180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="277" />
                    <RANKING place="1" resultid="2174" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26" number="42" gender="M" round="PRE" order="42">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="26000" number="0" />
                <HEAT heatid="26001" number="1" daytime="13:33" />
                <HEAT heatid="26002" number="2" daytime="13:34" />
                <HEAT heatid="26003" number="3" daytime="13:35" />
                <HEAT heatid="26004" number="4" daytime="13:36" />
                <HEAT heatid="26005" number="5" daytime="13:37" />
                <HEAT heatid="26006" number="6" daytime="13:38" />
                <HEAT heatid="26007" number="7" daytime="13:39" />
                <HEAT heatid="26008" number="8" daytime="13:40" />
                <HEAT heatid="26009" number="9" daytime="13:41" />
                <HEAT heatid="26010" number="10" daytime="13:41" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="5" resultid="139" />
                    <RANKING place="6" resultid="630" />
                    <RANKING place="3" resultid="1191" />
                    <RANKING place="7" resultid="1201" />
                    <RANKING place="1" resultid="1504" />
                    <RANKING place="9" resultid="1614" />
                    <RANKING place="4" resultid="1673" />
                    <RANKING place="2" resultid="1894" />
                    <RANKING place="8" resultid="2297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="9" resultid="108" />
                    <RANKING place="8" resultid="272" />
                    <RANKING place="3" resultid="517" />
                    <RANKING place="4" resultid="775" />
                    <RANKING place="2" resultid="1008" />
                    <RANKING place="7" resultid="1063" />
                    <RANKING place="1" resultid="1117" />
                    <RANKING place="10" resultid="1241" />
                    <RANKING place="5" resultid="1251" />
                    <RANKING place="12" resultid="1609" />
                    <RANKING place="11" resultid="1905" />
                    <RANKING place="6" resultid="2247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="4" resultid="390" />
                    <RANKING place="5" resultid="428" />
                    <RANKING place="3" resultid="448" />
                    <RANKING place="7" resultid="798" />
                    <RANKING place="1" resultid="950" />
                    <RANKING place="2" resultid="1097" />
                    <RANKING place="6" resultid="1330" />
                    <RANKING place="8" resultid="2022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="466" />
                    <RANKING place="2" resultid="846" />
                    <RANKING place="4" resultid="1365" />
                    <RANKING place="8" resultid="1418" />
                    <RANKING place="5" resultid="1473" />
                    <RANKING place="6" resultid="1523" />
                    <RANKING place="7" resultid="1595" />
                    <RANKING place="1" resultid="2151" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="45" number="43" gender="F" round="TIM" order="43">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="45000" number="0" />
                <HEAT heatid="45001" number="1" daytime="13:44" />
                <HEAT heatid="45002" number="2" daytime="13:46" />
                <HEAT heatid="45003" number="3" daytime="13:48" />
                <HEAT heatid="45004" number="4" daytime="13:50" />
                <HEAT heatid="45005" number="5" daytime="13:52" />
                <HEAT heatid="45006" number="6" daytime="13:54" />
                <HEAT heatid="45007" number="7" daytime="13:56" />
                <HEAT heatid="45008" number="8" daytime="13:58" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="60" />
                    <RANKING place="5" resultid="479" />
                    <RANKING place="3" resultid="1667" />
                    <RANKING place="6" resultid="2037" />
                    <RANKING place="4" resultid="2098" />
                    <RANKING place="1" resultid="2277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="170" />
                    <RANKING place="3" resultid="332" />
                    <RANKING place="5" resultid="641" />
                    <RANKING place="1" resultid="1247" />
                    <RANKING place="2" resultid="1979" />
                    <RANKING place="6" resultid="2187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="4" resultid="339" />
                    <RANKING place="5" resultid="624" />
                    <RANKING place="2" resultid="833" />
                    <RANKING place="1" resultid="1102" />
                    <RANKING place="3" resultid="1197" />
                    <RANKING place="8" resultid="1237" />
                    <RANKING place="7" resultid="1257" />
                    <RANKING place="6" resultid="1600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="791" />
                    <RANKING place="2" resultid="1134" />
                    <RANKING place="4" resultid="1575" />
                    <RANKING place="1" resultid="1709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="848" />
                    <RANKING place="2" resultid="1590" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="46" number="44" gender="M" round="TIM" order="44">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="46000" number="0" />
                <HEAT heatid="46001" number="1" daytime="14:02" />
                <HEAT heatid="46002" number="2" daytime="14:04" />
                <HEAT heatid="46003" number="3" daytime="14:06" />
                <HEAT heatid="46004" number="4" daytime="14:07" />
                <HEAT heatid="46005" number="5" daytime="14:09" />
                <HEAT heatid="46006" number="6" daytime="14:11" />
                <HEAT heatid="46007" number="7" daytime="14:12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="768" />
                    <RANKING place="2" resultid="1217" />
                    <RANKING place="3" resultid="1881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="10" resultid="84" />
                    <RANKING place="4" resultid="149" />
                    <RANKING place="11" resultid="175" />
                    <RANKING place="5" resultid="538" />
                    <RANKING place="7" resultid="654" />
                    <RANKING place="6" resultid="942" />
                    <RANKING place="3" resultid="946" />
                    <RANKING place="2" resultid="972" />
                    <RANKING place="1" resultid="1120" />
                    <RANKING place="12" resultid="1906" />
                    <RANKING place="9" resultid="1938" />
                    <RANKING place="8" resultid="2103" />
                    <RANKING place="13" resultid="2209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="4" resultid="87" />
                    <RANKING place="2" resultid="391" />
                    <RANKING place="1" resultid="429" />
                    <RANKING place="6" resultid="825" />
                    <RANKING place="3" resultid="841" />
                    <RANKING place="5" resultid="2023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="657" />
                    <RANKING place="1" resultid="809" />
                    <RANKING place="2" resultid="1474" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="31" number="45" gender="F" round="TIM" order="45">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="31000" number="0" />
                <HEAT heatid="31001" number="1" daytime="14:16" />
                <HEAT heatid="31002" number="2" daytime="14:18" />
                <HEAT heatid="31003" number="3" daytime="14:20" />
                <HEAT heatid="31004" number="4" daytime="14:21" />
                <HEAT heatid="31005" number="5" daytime="14:23" />
                <HEAT heatid="31006" number="6" daytime="14:25" />
                <HEAT heatid="31007" number="7" daytime="14:26" />
                <HEAT heatid="31008" number="8" daytime="14:28" />
                <HEAT heatid="31009" number="9" daytime="14:29" />
                <HEAT heatid="31010" number="10" daytime="14:31" />
                <HEAT heatid="31011" number="11" daytime="14:32" />
                <HEAT heatid="31012" number="12" daytime="14:34" />
                <HEAT heatid="31013" number="13" daytime="14:35" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="8" resultid="67" />
                    <RANKING place="4" resultid="227" />
                    <RANKING place="1" resultid="364" />
                    <RANKING place="7" resultid="480" />
                    <RANKING place="5" resultid="1668" />
                    <RANKING place="2" resultid="1740" />
                    <RANKING place="3" resultid="1802" />
                    <RANKING place="9" resultid="2038" />
                    <RANKING place="6" resultid="2099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="8" resultid="101" />
                    <RANKING place="4" resultid="125" />
                    <RANKING place="7" resultid="171" />
                    <RANKING place="1" resultid="333" />
                    <RANKING place="5" resultid="492" />
                    <RANKING place="9" resultid="642" />
                    <RANKING place="2" resultid="772" />
                    <RANKING place="6" resultid="1563" />
                    <RANKING place="3" resultid="2092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="14" resultid="144" />
                    <RANKING place="16" resultid="161" />
                    <RANKING place="13" resultid="340" />
                    <RANKING place="2" resultid="383" />
                    <RANKING place="10" resultid="416" />
                    <RANKING place="19" resultid="616" />
                    <RANKING place="4" resultid="620" />
                    <RANKING place="12" resultid="625" />
                    <RANKING place="6" resultid="649" />
                    <RANKING place="7" resultid="783" />
                    <RANKING place="1" resultid="1126" />
                    <RANKING place="9" resultid="1207" />
                    <RANKING place="15" resultid="1227" />
                    <RANKING place="3" resultid="1267" />
                    <RANKING place="8" resultid="1454" />
                    <RANKING place="17" resultid="1601" />
                    <RANKING place="5" resultid="1843" />
                    <RANKING place="11" resultid="1951" />
                    <RANKING place="18" resultid="2058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="4" resultid="157" />
                    <RANKING place="2" resultid="820" />
                    <RANKING place="3" resultid="1358" />
                    <RANKING place="6" resultid="1576" />
                    <RANKING place="1" resultid="1710" />
                    <RANKING place="5" resultid="2181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="278" />
                    <RANKING place="3" resultid="1508" />
                    <RANKING place="1" resultid="2175" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="32" number="46" gender="M" round="TIM" order="46">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <FEE value="700" currency="EUR" />
              <HEATS>
                <HEAT heatid="32000" number="0" />
                <HEAT heatid="32001" number="1" daytime="14:39" />
                <HEAT heatid="32002" number="2" daytime="14:41" />
                <HEAT heatid="32003" number="3" daytime="14:42" />
                <HEAT heatid="32004" number="4" daytime="14:44" />
                <HEAT heatid="32005" number="5" daytime="14:45" />
                <HEAT heatid="32006" number="6" daytime="14:47" />
                <HEAT heatid="32007" number="7" daytime="14:48" />
                <HEAT heatid="32008" number="8" daytime="14:49" />
                <HEAT heatid="32009" number="9" daytime="14:51" />
                <HEAT heatid="32010" number="10" daytime="14:52" />
                <HEAT heatid="32011" number="11" daytime="14:54" />
                <HEAT heatid="32012" number="12" daytime="14:55" />
                <HEAT heatid="32013" number="13" daytime="14:56" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="9" resultid="122" />
                    <RANKING place="10" resultid="177" />
                    <RANKING place="3" resultid="664" />
                    <RANKING place="5" resultid="1192" />
                    <RANKING place="8" resultid="1202" />
                    <RANKING place="7" resultid="1277" />
                    <RANKING place="6" resultid="1505" />
                    <RANKING place="2" resultid="1674" />
                    <RANKING place="4" resultid="1895" />
                    <RANKING place="1" resultid="2287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="6" resultid="63" />
                    <RANKING place="4" resultid="135" />
                    <RANKING place="3" resultid="150" />
                    <RANKING place="19" resultid="176" />
                    <RANKING place="13" resultid="273" />
                    <RANKING place="12" resultid="497" />
                    <RANKING place="10" resultid="776" />
                    <RANKING place="9" resultid="787" />
                    <RANKING place="7" resultid="813" />
                    <RANKING place="15" resultid="817" />
                    <RANKING place="1" resultid="1139" />
                    <RANKING place="18" resultid="1242" />
                    <RANKING place="11" resultid="1252" />
                    <RANKING place="16" resultid="1350" />
                    <RANKING place="21" resultid="1610" />
                    <RANKING place="5" resultid="1691" />
                    <RANKING place="2" resultid="1726" />
                    <RANKING place="8" resultid="1747" />
                    <RANKING place="23" resultid="1907" />
                    <RANKING place="20" resultid="1939" />
                    <RANKING place="17" resultid="2104" />
                    <RANKING place="22" resultid="2210" />
                    <RANKING place="14" resultid="2248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="2" resultid="392" />
                    <RANKING place="4" resultid="430" />
                    <RANKING place="3" resultid="449" />
                    <RANKING place="5" resultid="779" />
                    <RANKING place="6" resultid="799" />
                    <RANKING place="7" resultid="826" />
                    <RANKING place="1" resultid="1098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="467" />
                    <RANKING place="7" resultid="643" />
                    <RANKING place="8" resultid="683" />
                    <RANKING place="2" resultid="806" />
                    <RANKING place="3" resultid="1366" />
                    <RANKING place="6" resultid="1419" />
                    <RANKING place="4" resultid="1459" />
                    <RANKING place="5" resultid="1524" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="49" number="47" gender="F" round="TIM" order="47">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="49001" number="1" daytime="15:00" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="128" />
                    <RANKING place="2" resultid="1044" />
                    <RANKING place="1" resultid="1135" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="50" number="48" gender="M" round="TIM" order="48">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="50000" number="0" />
                <HEAT heatid="50001" number="1" daytime="15:03" />
                <HEAT heatid="50002" number="2" daytime="15:08" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="136" />
                    <RANKING place="1" resultid="1129" />
                    <RANKING place="3" resultid="1692" />
                    <RANKING place="4" resultid="1727" />
                    <RANKING place="5" resultid="2222" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="35" number="49" gender="F" round="TIM" order="49">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="35001" number="1" daytime="15:10" />
                <HEAT heatid="35002" number="2" daytime="15:14" />
                <HEAT heatid="35003" number="3" daytime="15:17" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="677" />
                    <RANKING place="2" resultid="1045" />
                    <RANKING place="1" resultid="1112" />
                    <RANKING place="5" resultid="1359" />
                    <RANKING place="4" resultid="1455" />
                    <RANKING place="6" resultid="1741" />
                    <RANKING place="3" resultid="1803" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="36" number="50" gender="M" round="TIM" order="50">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="36000" number="0" />
                <HEAT heatid="36001" number="1" daytime="15:23" />
                <HEAT heatid="36002" number="2" daytime="15:27" />
                <HEAT heatid="36003" number="3" daytime="15:30" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="518" />
                    <RANKING place="7" resultid="827" />
                    <RANKING place="1" resultid="951" />
                    <RANKING place="3" resultid="1009" />
                    <RANKING place="2" resultid="1367" />
                    <RANKING place="4" resultid="1596" />
                    <RANKING place="9" resultid="1875" />
                    <RANKING place="8" resultid="2071" />
                    <RANKING place="6" resultid="2288" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="53" number="51" gender="F" round="TIM" order="51">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="53000" number="0" />
                <HEAT heatid="53001" number="1" daytime="15:34" />
                <HEAT heatid="53002" number="2" daytime="15:38" />
                <HEAT heatid="53003" number="3" daytime="15:41" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="365" />
                    <RANKING place="2" resultid="2278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="1980" />
                    <RANKING place="2" resultid="2093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="3" resultid="384" />
                    <RANKING place="1" resultid="524" />
                    <RANKING place="2" resultid="1844" />
                    <RANKING place="4" resultid="1952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="2" resultid="792" />
                    <RANKING place="1" resultid="1711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="1509" />
                    <RANKING place="2" resultid="1591" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="54" number="52" gender="M" round="TIM" order="52">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="54001" number="1" daytime="15:44" />
                <HEAT heatid="54002" number="2" daytime="15:48" />
                <HEAT heatid="54003" number="3" daytime="15:51" />
                <HEAT heatid="54004" number="4" daytime="15:54" />
                <HEAT heatid="54005" number="5" daytime="15:57" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="1882" />
                    <RANKING place="1" resultid="1896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2009/2010">
                  <RANKINGS>
                    <RANKING place="7" resultid="498" />
                    <RANKING place="5" resultid="539" />
                    <RANKING place="6" resultid="943" />
                    <RANKING place="4" resultid="947" />
                    <RANKING place="2" resultid="973" />
                    <RANKING place="1" resultid="1121" />
                    <RANKING place="3" resultid="1130" />
                    <RANKING place="8" resultid="1351" />
                    <RANKING place="10" resultid="1940" />
                    <RANKING place="9" resultid="2249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="2" resultid="450" />
                    <RANKING place="3" resultid="842" />
                    <RANKING place="1" resultid="952" />
                    <RANKING place="4" resultid="2024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2006 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="1159" />
                    <RANKING place="1" resultid="1368" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="55" number="141" gender="F" round="FIN" order="53">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="55001" number="1" daytime="16:30" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="2347" />
                    <RANKING place="7" resultid="2348" />
                    <RANKING place="6" resultid="2349" />
                    <RANKING place="8" resultid="2350" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="56" number="241" gender="F" round="FIN" order="54">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="56001" number="1" daytime="16:32" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="13" name="2012 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2351" />
                    <RANKING place="2" resultid="2352" />
                    <RANKING place="3" resultid="2353" />
                    <RANKING place="4" resultid="2354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2351" />
                    <RANKING place="2" resultid="2352" />
                    <RANKING place="3" resultid="2353" />
                    <RANKING place="4" resultid="2354" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="57" number="142" gender="M" round="FIN" order="55">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="57001" number="1" daytime="16:35" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2355" />
                    <RANKING place="2" resultid="2356" />
                    <RANKING place="3" resultid="2357" />
                    <RANKING place="4" resultid="2358" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="58" number="242" gender="M" round="FIN" order="56">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="58001" number="1" daytime="16:38" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="14" name="2011 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2359" />
                    <RANKING place="2" resultid="2360" />
                    <RANKING place="3" resultid="2361" />
                    <RANKING place="4" resultid="2362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Juniorenwertung" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="59" number="125" gender="F" round="FIN" order="57">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="59001" number="1" daytime="16:54" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="2315" />
                    <RANKING place="3" resultid="2316" />
                    <RANKING place="5" resultid="2317" />
                    <RANKING place="6" resultid="2318" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="60" number="225" gender="F" round="FIN" order="58">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="60001" number="1" daytime="16:57" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="13" name="2012 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2319" />
                    <RANKING place="2" resultid="2320" />
                    <RANKING place="3" resultid="2321" />
                    <RANKING place="4" resultid="2322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2320" />
                    <RANKING place="2" resultid="2322" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="61" number="126" gender="M" round="FIN" order="59">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="61001" number="1" daytime="17:00" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="2323" />
                    <RANKING place="5" resultid="2324" />
                    <RANKING place="4" resultid="2325" />
                    <RANKING place="6" resultid="2326" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="62" number="226" gender="M" round="FIN" order="60">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="62001" number="1" daytime="17:03" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="14" name="2011 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2327" />
                    <RANKING place="2" resultid="2328" />
                    <RANKING place="3" resultid="2329" />
                    <RANKING place="4" resultid="2330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2328" />
                    <RANKING place="2" resultid="2329" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="63" number="139" gender="F" round="FIN" order="61">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="63001" number="1" daytime="17:19" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="2331" />
                    <RANKING place="6" resultid="2332" />
                    <RANKING place="5" resultid="2333" />
                    <RANKING place="7" resultid="2334" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="64" number="239" gender="F" round="FIN" order="62">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="64001" number="1" daytime="17:22" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="13" name="2012 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2335" />
                    <RANKING place="3" resultid="2336" />
                    <RANKING place="2" resultid="2337" />
                    <RANKING place="4" resultid="2338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2335" />
                    <RANKING place="2" resultid="2336" />
                    <RANKING place="3" resultid="2338" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="65" number="140" gender="M" round="FIN" order="63">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="65001" number="1" daytime="17:25" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="2339" />
                    <RANKING place="4" resultid="2340" />
                    <RANKING place="3" resultid="2341" />
                    <RANKING place="5" resultid="2342" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="66" number="240" gender="M" round="FIN" order="64">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="66001" number="1" daytime="17:27" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="14" name="2011 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2343" />
                    <RANKING place="2" resultid="2344" />
                    <RANKING place="4" resultid="2345" />
                    <RANKING place="3" resultid="2346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2345" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="67" number="123" gender="F" round="FIN" order="65">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="67000" number="0" />
                <HEAT heatid="67001" number="1" daytime="17:43" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="2299" />
                    <RANKING place="7" resultid="2300" />
                    <RANKING place="6" resultid="2301" />
                    <RANKING place="8" resultid="2302" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="68" number="223" gender="F" round="FIN" order="66">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="68001" number="1" daytime="17:46" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="13" name="2012 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2303" />
                    <RANKING place="2" resultid="2304" />
                    <RANKING place="3" resultid="2305" />
                    <RANKING place="4" resultid="2306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2303" />
                    <RANKING place="2" resultid="2304" />
                    <RANKING place="3" resultid="2305" />
                    <RANKING place="4" resultid="2306" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="69" number="124" gender="M" round="FIN" order="67">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="69001" number="1" daytime="17:49" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="17" agemin="12" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="2307" />
                    <RANKING place="1" resultid="2308" />
                    <RANKING place="3" resultid="2309" />
                    <RANKING place="2" resultid="2310" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="70" number="224" gender="M" round="FIN" order="68">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="70001" number="1" daytime="17:52" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="14" name="2011 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2311" />
                    <RANKING place="4" resultid="2312" />
                    <RANKING place="2" resultid="2313" />
                    <RANKING place="3" resultid="2314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Juniorenwertung" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="71" number="53" gender="F" round="TIM" order="69">
              <SWIMSTYLE stroke="MEDLEY" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="71001" number="1" daytime="18:07" />
                <HEAT heatid="71002" number="2" daytime="18:10" />
                <HEAT heatid="71003" number="3" daytime="18:13" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Jahrgänge 2015 und älter">
                  <RANKINGS>
                    <RANKING place="5" resultid="283" />
                    <RANKING place="7" resultid="609" />
                    <RANKING place="4" resultid="765" />
                    <RANKING place="1" resultid="851" />
                    <RANKING place="2" resultid="1179" />
                    <RANKING place="3" resultid="1286" />
                    <RANKING place="6" resultid="1848" />
                    <RANKING place="8" resultid="1854" />
                    <RANKING place="9" resultid="1860" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="72" number="54" gender="M" round="TIM" order="70">
              <SWIMSTYLE stroke="MEDLEY" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="72001" number="1" daytime="18:18" />
                <HEAT heatid="72002" number="2" daytime="18:21" />
                <HEAT heatid="72003" number="3" daytime="18:23" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Jahrgänge 2015 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="284" />
                    <RANKING place="7" resultid="607" />
                    <RANKING place="4" resultid="763" />
                    <RANKING place="2" resultid="852" />
                    <RANKING place="5" resultid="853" />
                    <RANKING place="8" resultid="854" />
                    <RANKING place="9" resultid="1181" />
                    <RANKING place="3" resultid="1284" />
                    <RANKING place="6" resultid="1846" />
                    <RANKING place="10" resultid="1852" />
                    <RANKING place="11" resultid="1858" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="ATSV Freiberg e.V." nation="GER" region="12" code="3324">
          <ATHLETES>
            <ATHLETE athleteid="50" birthdate="2013-01-01" gender="M" lastname="Ahlbrecht" firstname="Theo" license="484744" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:38.75" heatid="4015" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:31.27" heatid="8024" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:24.39" heatid="10012" lane="4" />
                <ENTRY eventid="14" entrytime="00:00:38.10" heatid="14007" lane="4" />
                <ENTRY eventid="16" entrytime="00:01:23.46" heatid="16010" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:09.82" heatid="20021" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="181" eventid="4" swimtime="00:00:38.01" lane="1" heatid="4015" points="196" />
                <RESULT resultid="182" eventid="8" swimtime="00:00:31.47" lane="4" heatid="8024" points="262" />
                <RESULT resultid="183" eventid="10" swimtime="00:01:23.05" lane="4" heatid="10012" points="208">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="184" eventid="14" swimtime="00:00:38.05" lane="4" heatid="14007" points="186" />
                <RESULT resultid="185" eventid="16" swimtime="00:01:22.70" lane="2" heatid="16010" points="199">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="186" eventid="20" swimtime="00:01:10.67" lane="3" heatid="20021" points="255">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="51" birthdate="2013-01-01" gender="F" lastname="Brocke" firstname="Fiene" license="445947" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:43.85" heatid="3016" lane="4" />
                <ENTRY eventid="5" entrytime="00:01:43.57" heatid="5009" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:38.09" heatid="7018" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:47.52" heatid="13006" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:47.83" heatid="17013" lane="1" />
                <ENTRY eventid="21" entrytime="00:03:21.71" heatid="21002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="187" eventid="3" swimtime="00:00:42.61" lane="4" heatid="3016" points="208" />
                <RESULT resultid="188" eventid="5" swimtime="00:01:42.69" lane="1" heatid="5009" points="223">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="189" eventid="7" swimtime="00:00:36.97" lane="2" heatid="7018" points="238" />
                <RESULT resultid="190" eventid="13" swimtime="00:00:42.05" lane="3" heatid="13006" points="194" />
                <RESULT resultid="191" eventid="17" swimtime="00:00:47.34" lane="1" heatid="17013" points="215" />
                <RESULT resultid="192" eventid="21" swimtime="00:03:17.30" lane="1" heatid="21002" points="235">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                    <SPLIT distance="100" swimtime="00:01:35.03" />
                    <SPLIT distance="150" swimtime="00:02:31.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="52" birthdate="2014-01-01" gender="F" lastname="Ferkinghoff" firstname="Helene" license="445062" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:41.02" heatid="3018" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:34.10" heatid="7025" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:37.02" heatid="9007" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:42.31" heatid="13009" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:30.03" heatid="15013" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:19.49" heatid="19020" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="193" eventid="3" swimtime="00:00:40.06" lane="4" heatid="3018" points="250" />
                <RESULT resultid="194" eventid="7" swimtime="00:00:34.22" lane="3" heatid="7025" points="300" />
                <RESULT resultid="195" eventid="9" swimtime="00:01:31.77" lane="2" heatid="9007" points="233">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="196" eventid="13" swimtime="00:00:41.63" lane="2" heatid="13009" points="200" />
                <RESULT resultid="197" eventid="15" swimtime="00:01:31.92" lane="4" heatid="15013" points="212">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="198" eventid="19" swimtime="00:01:19.57" lane="1" heatid="19020" points="251">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="53" birthdate="2014-01-01" gender="F" lastname="Grämer" firstname="Stella" license="445949" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:39.59" heatid="3022" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:34.94" heatid="7024" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:27.66" heatid="9012" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:37.99" heatid="13011" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:24.44" heatid="15014" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:19.69" heatid="19019" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="199" eventid="3" swimtime="00:00:39.28" lane="4" heatid="3022" points="265" />
                <RESULT resultid="200" eventid="7" swimtime="00:00:34.43" lane="1" heatid="7024" points="295" />
                <RESULT resultid="201" eventid="9" swimtime="00:01:31.22" lane="2" heatid="9012" points="237">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="202" eventid="13" swimtime="00:00:39.91" lane="3" heatid="13011" points="227" />
                <RESULT resultid="203" eventid="15" swimtime="00:01:31.16" lane="1" heatid="15014" points="218">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="204" eventid="19" swimtime="00:01:21.57" lane="2" heatid="19019" points="233">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="54" birthdate="2015-01-01" gender="F" lastname="Heinz" firstname="Elizabeth" license="471931" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:40.86" heatid="3021" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:36.61" heatid="7021" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:35.62" heatid="9009" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:43.29" heatid="13014" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:29.56" heatid="15013" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:46.77" heatid="17018" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="205" eventid="3" swimtime="00:00:40.89" lane="3" heatid="3021" points="235" />
                <RESULT resultid="206" eventid="7" swimtime="00:00:35.46" lane="1" heatid="7021" points="270" />
                <RESULT resultid="207" eventid="9" swimtime="00:01:32.28" lane="3" heatid="9009" points="229">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="208" eventid="13" swimtime="00:00:42.80" lane="4" heatid="13014" points="184" />
                <RESULT resultid="209" eventid="15" swimtime="00:01:31.28" lane="1" heatid="15013" points="217">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="210" eventid="17" swimtime="00:00:48.38" lane="4" heatid="17018" points="201" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="55" birthdate="2014-01-01" gender="F" lastname="Irmscher" firstname="Nora" license="445948" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:44.43" heatid="1002" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:35.46" heatid="7023" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:37.53" heatid="9007" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:43.87" heatid="13008" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:51.67" heatid="17010" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:23.86" heatid="19016" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="211" eventid="1" swimtime="00:01:46.42" lane="1" heatid="1002" points="131">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="212" eventid="7" swimtime="00:00:36.04" lane="2" heatid="7023" points="257" />
                <RESULT resultid="213" eventid="9" swimtime="00:01:37.44" lane="3" heatid="9007" points="195">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="214" eventid="13" swimtime="00:00:44.83" lane="3" heatid="13008" points="160" />
                <RESULT resultid="215" eventid="17" swimtime="00:00:51.73" lane="4" heatid="17010" points="164" />
                <RESULT resultid="216" eventid="19" swimtime="00:01:22.19" lane="1" heatid="19016" points="228">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="56" birthdate="2016-01-01" gender="M" lastname="Kaiser" firstname="Tom" license="476731" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:55.17" heatid="4002" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:44.04" heatid="8006" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:53.15" heatid="10002" lane="1" />
                <ENTRY eventid="14" entrytime="00:01:13.61" heatid="14001" lane="3" />
                <ENTRY eventid="18" entrytime="00:01:00.43" heatid="18002" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:40.44" heatid="20004" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="217" eventid="4" swimtime="00:00:55.34" lane="3" heatid="4002" points="63" />
                <RESULT resultid="218" eventid="8" swimtime="00:00:44.46" lane="2" heatid="8006" points="93" />
                <RESULT resultid="219" eventid="10" swimtime="00:02:00.95" lane="1" heatid="10002" points="67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="220" eventid="14" status="DNS" swimtime="00:00:00.00" lane="3" heatid="14001" />
                <RESULT resultid="221" eventid="18" swimtime="00:00:58.66" lane="3" heatid="18002" points="76" />
                <RESULT resultid="222" eventid="20" swimtime="00:01:39.96" lane="3" heatid="20004" points="90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="57" birthdate="2012-01-01" gender="F" lastname="Kaiser" firstname="Zoe" license="431997" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.24" heatid="43010" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:46.74" heatid="27002" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:33.14" heatid="41008" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:35.74" heatid="25005" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:09.36" heatid="31009" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="223" eventid="43" swimtime="00:00:30.34" lane="1" heatid="43010" points="431" />
                <RESULT resultid="224" eventid="27" swimtime="00:00:46.93" lane="4" heatid="27002" points="220" />
                <RESULT resultid="225" eventid="41" swimtime="00:00:34.55" lane="3" heatid="41008" points="351" />
                <RESULT resultid="226" eventid="25" swimtime="00:00:36.09" lane="1" heatid="25005" points="342" />
                <RESULT resultid="227" eventid="31" swimtime="00:01:11.53" lane="3" heatid="31009" points="346">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="58" birthdate="2015-01-01" gender="M" lastname="Kononchuk" firstname="Georgii" license="500287" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:49.34" heatid="4006" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:40.82" heatid="8010" lane="4" />
                <ENTRY eventid="10" entrytime="00:00:00.00" heatid="10001" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:49.86" heatid="16008" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:34.22" heatid="20007" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="228" eventid="4" swimtime="00:00:51.49" lane="3" heatid="4006" points="79" />
                <RESULT resultid="229" eventid="8" swimtime="00:00:43.01" lane="4" heatid="8010" points="102" />
                <RESULT resultid="230" eventid="10" status="DSQ" swimtime="00:01:52.79" lane="3" heatid="10001" comment="Die Arme wurden während der Schwimmstrecke nicht gleichzeitig über Wasser nach vorn gebracht.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="231" eventid="16" swimtime="00:02:01.01" lane="4" heatid="16008" points="63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="232" eventid="20" swimtime="00:01:45.17" lane="2" heatid="20007" points="77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="59" birthdate="2013-01-01" gender="M" lastname="Oehme" firstname="Arvid" license="445060" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:20.86" heatid="2005" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:31.63" heatid="8019" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:23.59" heatid="10012" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:34.05" heatid="14011" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:44.20" heatid="18008" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:12.89" heatid="20016" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="233" eventid="2" status="DNS" swimtime="00:00:00.00" lane="2" heatid="2005" />
                <RESULT resultid="234" eventid="8" status="DNS" swimtime="00:00:00.00" lane="2" heatid="8019" />
                <RESULT resultid="235" eventid="10" status="DNS" swimtime="00:00:00.00" lane="1" heatid="10012" />
                <RESULT resultid="236" eventid="14" status="DNS" swimtime="00:00:00.00" lane="3" heatid="14011" />
                <RESULT resultid="237" eventid="18" status="DNS" swimtime="00:00:00.00" lane="2" heatid="18008" />
                <RESULT resultid="238" eventid="20" status="DNS" swimtime="00:00:00.00" lane="1" heatid="20016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="60" birthdate="2016-01-01" gender="F" lastname="Paech" firstname="Eveline" license="500288" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:57.89" heatid="3005" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:47.27" heatid="7009" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:53.80" heatid="15005" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:00.00" heatid="17001" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:44.74" heatid="19007" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="239" eventid="3" swimtime="00:00:53.19" lane="1" heatid="3005" points="106" />
                <RESULT resultid="240" eventid="7" swimtime="00:00:42.93" lane="3" heatid="7009" points="152" />
                <RESULT resultid="241" eventid="15" swimtime="00:02:10.17" lane="2" heatid="15005" points="74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="242" eventid="17" swimtime="00:01:08.46" lane="3" heatid="17001" points="71" />
                <RESULT resultid="243" eventid="19" swimtime="00:01:58.71" lane="4" heatid="19007" points="75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="61" birthdate="2013-01-01" gender="F" lastname="Queck" firstname="Fabienne" license="451852" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:40.01" heatid="3018" lane="2" />
                <ENTRY eventid="5" entrytime="00:01:33.48" heatid="5015" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:31.08" heatid="9011" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:41.57" heatid="13010" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:28.86" heatid="15013" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:41.24" heatid="17020" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="244" eventid="3" swimtime="00:00:39.44" lane="2" heatid="3018" points="262" />
                <RESULT resultid="245" eventid="5" swimtime="00:01:31.51" lane="3" heatid="5015" points="316">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="246" eventid="9" swimtime="00:01:28.22" lane="3" heatid="9011" points="262">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="247" eventid="13" swimtime="00:00:40.84" lane="4" heatid="13010" points="212" />
                <RESULT resultid="248" eventid="15" swimtime="00:01:30.76" lane="3" heatid="15013" points="221">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="249" eventid="17" swimtime="00:00:42.32" lane="3" heatid="17020" points="301" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="62" birthdate="2014-01-01" gender="F" lastname="Riedel" firstname="Hely Margo" license="445061" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:22.08" heatid="1004" lane="2" />
                <ENTRY eventid="5" entrytime="00:01:23.94" heatid="5014" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:30.84" heatid="7029" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:33.99" heatid="13015" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:18.62" heatid="15018" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:09.72" heatid="19024" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="250" eventid="1" swimtime="00:01:18.59" lane="2" heatid="1004" points="325">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="251" eventid="5" swimtime="00:01:27.17" lane="2" heatid="5014" points="366">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="252" eventid="7" swimtime="00:00:31.30" lane="2" heatid="7029" points="393" />
                <RESULT resultid="253" eventid="13" swimtime="00:00:34.30" lane="2" heatid="13015" points="359" />
                <RESULT resultid="254" eventid="15" swimtime="00:01:18.60" lane="3" heatid="15018" points="340">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="255" eventid="19" swimtime="00:01:10.62" lane="2" heatid="19024" points="360">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="63" birthdate="2011-01-01" gender="M" lastname="Rülke" firstname="Luca" license="431995" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:34.11" heatid="44001" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:43.73" heatid="28001" lane="2" />
                <ENTRY eventid="48" entrytime="00:01:27.03" heatid="48001" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:42.31" heatid="42001" lane="1" />
                <ENTRY eventid="26" entrytime="00:00:44.32" heatid="26001" lane="3" />
                <ENTRY eventid="32" entrytime="00:01:15.33" heatid="32002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="256" eventid="44" swimtime="00:00:33.17" lane="2" heatid="44001" points="224" />
                <RESULT resultid="257" eventid="28" swimtime="00:00:43.79" lane="2" heatid="28001" points="184" />
                <RESULT resultid="258" eventid="48" swimtime="00:01:30.51" lane="1" heatid="48001" points="152">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="259" eventid="42" status="DNS" swimtime="00:00:00.00" lane="1" heatid="42001" />
                <RESULT resultid="260" eventid="26" status="DNS" swimtime="00:00:00.00" lane="3" heatid="26001" />
                <RESULT resultid="261" eventid="32" status="DNS" swimtime="00:00:00.00" lane="4" heatid="32002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="64" birthdate="2012-01-01" gender="M" lastname="Tanneberger" firstname="Arian" license="434981" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:19.72" heatid="2006" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:29.44" heatid="8025" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:18.17" heatid="10013" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:34.33" heatid="14012" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:38.17" heatid="18015" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:07.87" heatid="20022" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="262" eventid="2" swimtime="00:01:18.20" lane="1" heatid="2006" points="228">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="263" eventid="8" swimtime="00:00:29.65" lane="3" heatid="8025" points="314" />
                <RESULT resultid="264" eventid="10" swimtime="00:01:16.49" lane="3" heatid="10013" points="267">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="265" eventid="14" swimtime="00:00:34.39" lane="1" heatid="14012" points="252" />
                <RESULT resultid="266" eventid="18" swimtime="00:00:37.73" lane="4" heatid="18015" points="289" />
                <RESULT resultid="267" eventid="20" swimtime="00:01:06.95" lane="4" heatid="20022" points="300">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="65" birthdate="2010-01-01" gender="M" lastname="Tanneberger" firstname="Janis" license="407515" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.45" heatid="44009" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:34.96" heatid="28005" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:10.62" heatid="34005" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:30.72" heatid="42004" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:33.15" heatid="26004" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:02.26" heatid="32006" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="268" eventid="44" swimtime="00:00:27.44" lane="4" heatid="44009" points="396" />
                <RESULT resultid="269" eventid="28" swimtime="00:00:35.75" lane="1" heatid="28005" points="339" />
                <RESULT resultid="270" eventid="34" swimtime="00:01:12.00" lane="4" heatid="34005" points="320">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="271" eventid="42" swimtime="00:00:30.77" lane="3" heatid="42004" points="353" />
                <RESULT resultid="272" eventid="26" swimtime="00:00:33.26" lane="1" heatid="26004" points="293" />
                <RESULT resultid="273" eventid="32" swimtime="00:01:03.41" lane="4" heatid="32006" points="353">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="66" birthdate="2003-01-01" gender="F" lastname="Wolf" firstname="Leonie" license="242026" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:29.26" heatid="43014" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:15.78" heatid="33010" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:32.28" heatid="41012" lane="4" />
                <ENTRY eventid="25" entrytime="00:00:34.05" heatid="25009" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:06.15" heatid="31013" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="274" eventid="43" swimtime="00:00:29.97" lane="3" heatid="43014" points="447" />
                <RESULT resultid="275" eventid="33" swimtime="00:01:17.95" lane="3" heatid="33010" points="381">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="276" eventid="41" swimtime="00:00:33.62" lane="4" heatid="41012" points="381" />
                <RESULT resultid="277" eventid="25" swimtime="00:00:34.83" lane="3" heatid="25009" points="380" />
                <RESULT resultid="278" eventid="31" swimtime="00:01:08.14" lane="3" heatid="31013" points="401">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:14.15" lane="1" heatid="11002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="178" eventid="11" swimtime="00:02:36.61" lane="1" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:09.41" />
                    <SPLIT distance="150" swimtime="00:01:54.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="53" number="1" />
                    <RELAYPOSITION athleteid="55" number="2" />
                    <RELAYPOSITION athleteid="58" number="3" />
                    <RELAYPOSITION athleteid="56" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:13.30" lane="3" heatid="11002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="179" eventid="11" swimtime="00:02:05.42" lane="3" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:04.15" />
                    <SPLIT distance="150" swimtime="00:01:35.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="64" number="1" />
                    <RELAYPOSITION athleteid="52" number="2" />
                    <RELAYPOSITION athleteid="50" number="3" />
                    <RELAYPOSITION athleteid="62" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="23" entrytime="00:02:20.00" lane="3" heatid="23003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="180" eventid="23" swimtime="00:02:22.37" lane="3" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:17.32" />
                    <SPLIT distance="150" swimtime="00:01:51.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="62" number="1" />
                    <RELAYPOSITION athleteid="61" number="2" />
                    <RELAYPOSITION athleteid="64" number="3" />
                    <RELAYPOSITION athleteid="50" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Dresdner Delphine e.V." nation="GER" region="12" code="5753">
          <ATHLETES>
            <ATHLETE athleteid="1" birthdate="2016-01-01" gender="M" lastname="Asanow" firstname="Michael" license="463183" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:44.16" heatid="4012" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:38.70" heatid="8021" lane="1" />
                <ENTRY eventid="14" entrytime="00:01:00.00" heatid="14002" lane="1" />
                <ENTRY eventid="16" entrytime="00:01:40.00" heatid="16007" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:33.36" heatid="20018" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1" eventid="4" swimtime="00:00:45.39" lane="2" heatid="4012" points="115" />
                <RESULT resultid="2" eventid="8" swimtime="00:00:38.55" lane="1" heatid="8021" points="143" />
                <RESULT resultid="3" eventid="14" swimtime="00:00:48.49" lane="1" heatid="14002" points="90" />
                <RESULT resultid="4" eventid="16" swimtime="00:01:35.25" lane="3" heatid="16007" points="130">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5" eventid="20" swimtime="00:01:25.76" lane="4" heatid="20018" points="142">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="2" birthdate="2013-01-01" gender="M" lastname="Barthel" firstname="Lennard" license="437409" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:31.60" heatid="2005" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:34.59" heatid="8016" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:27.43" heatid="10006" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:36.95" heatid="14007" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:13.69" heatid="20015" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="6" eventid="2" swimtime="00:01:18.07" lane="4" heatid="2005" points="229">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="7" eventid="8" swimtime="00:00:33.42" lane="3" heatid="8016" points="219" />
                <RESULT resultid="8" eventid="10" swimtime="00:01:22.19" lane="2" heatid="10006" points="215">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="9" eventid="14" swimtime="00:00:35.13" lane="2" heatid="14007" points="237" />
                <RESULT resultid="10" eventid="20" swimtime="00:01:13.51" lane="2" heatid="20015" points="226">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="3" birthdate="2016-01-01" gender="F" lastname="Böck" firstname="Merle" license="479066" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:46.89" heatid="3012" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:39.60" heatid="7017" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:50.00" heatid="15006" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:36.97" heatid="19010" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="11" eventid="3" swimtime="00:00:46.24" lane="2" heatid="3012" points="162" />
                <RESULT resultid="12" eventid="7" swimtime="00:00:38.25" lane="4" heatid="7017" points="215" />
                <RESULT resultid="13" eventid="15" swimtime="00:01:45.63" lane="2" heatid="15006" points="140">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="14" eventid="19" swimtime="00:01:39.29" lane="4" heatid="19010" points="129">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="4" birthdate="2016-01-01" gender="F" lastname="Göllner" firstname="Lisbeth" license="463213" nation="GER">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:00:36.12" heatid="7027" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:42.85" heatid="13013" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:45.59" heatid="15008" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:47.05" heatid="17017" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:28.11" heatid="19014" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="15" eventid="7" swimtime="00:00:36.53" lane="3" heatid="7027" points="247" />
                <RESULT resultid="16" eventid="13" swimtime="00:00:43.41" lane="3" heatid="13013" points="177" />
                <RESULT resultid="17" eventid="15" swimtime="00:01:36.30" lane="4" heatid="15008" points="185">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="18" eventid="17" swimtime="00:00:47.55" lane="2" heatid="17017" points="212" />
                <RESULT resultid="19" eventid="19" swimtime="00:01:27.82" lane="1" heatid="19014" points="187">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="5" birthdate="2016-01-01" gender="M" lastname="Graf" firstname="Theodor Alexander" license="463231" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:50.79" heatid="4005" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:46.52" heatid="8005" lane="3" />
                <ENTRY eventid="18" entrytime="00:01:05.21" heatid="18002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="20" eventid="4" swimtime="00:00:53.04" lane="1" heatid="4005" points="72" />
                <RESULT resultid="21" eventid="8" swimtime="00:00:46.06" lane="3" heatid="8005" points="83" />
                <RESULT resultid="22" eventid="18" swimtime="00:01:00.58" lane="4" heatid="18002" points="69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="6" birthdate="2016-01-01" gender="F" lastname="Herrmann" firstname="Caroline" license="480714" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:51.42" heatid="3009" lane="3" />
                <ENTRY eventid="5" entrytime="00:02:00.00" heatid="5003" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:44.45" heatid="7010" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:55.06" heatid="17006" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="23" eventid="3" status="DSQ" swimtime="00:00:51.77" lane="3" heatid="3009" comment="Die Sportlerin hat bei der Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt." />
                <RESULT resultid="24" eventid="5" swimtime="00:02:00.58" lane="2" heatid="5003" points="138">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="25" eventid="7" swimtime="00:00:44.25" lane="2" heatid="7010" points="139" />
                <RESULT resultid="26" eventid="17" swimtime="00:00:52.86" lane="2" heatid="17006" points="154" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="7" birthdate="2016-01-01" gender="F" lastname="Marr" firstname="Vanessa" license="479065" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:46.17" heatid="3000" lane="0" />
                <ENTRY eventid="5" entrytime="00:01:53.34" heatid="5000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:42.61" heatid="7000" lane="0" />
                <ENTRY eventid="15" entrytime="00:01:50.00" heatid="15000" lane="0" />
                <ENTRY eventid="17" entrytime="00:00:53.28" heatid="17000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="27" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="28" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="29" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="30" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="31" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="8" birthdate="2016-01-01" gender="M" lastname="Neumann" firstname="Philipp" license="463221" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:51.82" heatid="4004" lane="1" />
                <ENTRY eventid="6" entrytime="00:01:53.20" heatid="6008" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:43.48" heatid="8007" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:51.89" heatid="18011" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="32" eventid="4" swimtime="00:00:47.47" lane="1" heatid="4004" points="101" />
                <RESULT resultid="33" eventid="6" swimtime="00:01:49.30" lane="3" heatid="6008" points="129">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="34" eventid="8" swimtime="00:00:43.99" lane="4" heatid="8007" points="96" />
                <RESULT resultid="35" eventid="18" swimtime="00:00:49.93" lane="3" heatid="18011" points="124" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="9" birthdate="2016-01-01" gender="F" lastname="Pinera de la Cruz" firstname="Annabell" license="464581" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:46.99" heatid="3012" lane="3" />
                <ENTRY eventid="5" entrytime="00:01:52.36" heatid="5012" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:44.13" heatid="7011" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:53.11" heatid="17008" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="36" eventid="3" swimtime="00:00:48.46" lane="3" heatid="3012" points="141" />
                <RESULT resultid="37" eventid="5" swimtime="00:01:51.09" lane="4" heatid="5012" points="176">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="38" eventid="7" swimtime="00:00:43.22" lane="3" heatid="7011" points="149" />
                <RESULT resultid="39" eventid="17" swimtime="00:00:54.66" lane="2" heatid="17008" points="139" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="10" birthdate="2016-01-01" gender="F" lastname="Reichelt" firstname="Anna" license="463228" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:45.36" heatid="3020" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:36.07" heatid="7027" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:39.07" heatid="9015" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:46.16" heatid="13013" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:24.39" heatid="19022" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="40" eventid="3" swimtime="00:00:43.57" lane="4" heatid="3020" points="194" />
                <RESULT resultid="41" eventid="7" swimtime="00:00:35.01" lane="2" heatid="7027" points="280" />
                <RESULT resultid="42" eventid="9" swimtime="00:01:36.41" lane="2" heatid="9015" points="201">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="43" eventid="13" swimtime="00:00:46.39" lane="4" heatid="13013" points="145" />
                <RESULT resultid="44" eventid="19" swimtime="00:01:21.23" lane="3" heatid="19022" points="236">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="11" birthdate="2016-01-01" gender="F" lastname="Scale" firstname="Magdalena" license="485561" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:53.97" heatid="3006" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:47.61" heatid="7009" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:57.25" heatid="17006" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="45" eventid="3" swimtime="00:00:49.84" lane="2" heatid="3006" points="130" />
                <RESULT resultid="46" eventid="7" swimtime="00:00:44.34" lane="4" heatid="7009" points="138" />
                <RESULT resultid="47" eventid="17" swimtime="00:00:53.79" lane="4" heatid="17006" points="146" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="12" birthdate="2016-01-01" gender="F" lastname="Sendrowski" firstname="Lena Sophie" license="464953" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:58.99" heatid="5004" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:42.99" heatid="7012" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:56.30" heatid="13002" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:54.31" heatid="17008" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="48" eventid="5" swimtime="00:01:53.57" lane="4" heatid="5004" points="165">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="49" eventid="7" swimtime="00:00:42.39" lane="3" heatid="7012" points="158" />
                <RESULT resultid="50" eventid="13" swimtime="00:00:49.20" lane="3" heatid="13002" points="121" />
                <RESULT resultid="51" eventid="17" swimtime="00:00:53.44" lane="4" heatid="17008" points="149" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="13" birthdate="2016-01-01" gender="F" lastname="Wollmann" firstname="Maja" license="463178" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.73" heatid="3000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:40.56" heatid="7000" lane="0" />
                <ENTRY eventid="9" entrytime="00:01:38.33" heatid="9000" lane="0" />
                <ENTRY eventid="13" entrytime="00:00:47.30" heatid="13000" lane="0" />
                <ENTRY eventid="15" entrytime="00:01:35.75" heatid="15000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="52" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="53" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="54" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
                <RESULT resultid="55" eventid="13" status="WDR" swimtime="00:00:00.00" lane="0" heatid="13000" />
                <RESULT resultid="56" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="FC Erzgebirge Aue" nation="GER" region="12" code="7123">
          <ATHLETES>
            <ATHLETE athleteid="128" birthdate="2012-01-01" gender="M" lastname="Leonhardt" firstname="Jonas" license="482422" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:39.25" heatid="4016" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:32.15" heatid="8019" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:29.36" heatid="16011" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:14.50" heatid="20014" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="598" eventid="4" swimtime="00:00:37.60" lane="3" heatid="4016" points="203" />
                <RESULT resultid="599" eventid="8" swimtime="00:00:32.02" lane="3" heatid="8019" points="249" />
                <RESULT resultid="600" eventid="16" swimtime="00:01:26.92" lane="4" heatid="16011" points="171">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="601" eventid="20" swimtime="00:01:13.07" lane="2" heatid="20014" points="231">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129" birthdate="2012-01-01" gender="M" lastname="Weigel" firstname="Richard" license="482426" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:40.08" heatid="4016" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:34.83" heatid="8015" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:28.34" heatid="16011" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:46.48" heatid="18007" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="602" eventid="4" swimtime="00:00:42.97" lane="1" heatid="4016" points="136" />
                <RESULT resultid="603" eventid="8" swimtime="00:00:34.63" lane="3" heatid="8015" points="197" />
                <RESULT resultid="604" eventid="16" swimtime="00:01:30.72" lane="1" heatid="16011" points="151">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="605" eventid="18" swimtime="00:00:50.02" lane="2" heatid="18007" points="124" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Freibadverein Bad Blankenburg" nation="GER" region="16" code="7328">
          <ATHLETES>
            <ATHLETE athleteid="264" birthdate="2006-01-01" gender="M" lastname="Döring" firstname="Ferdinand" license="354729" nation="GER">
              <ENTRIES>
                <ENTRY eventid="30" entrytime="00:01:00.30" heatid="30006" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:03.12" heatid="34005" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:26.91" heatid="42008" lane="2" />
                <ENTRY eventid="54" entrytime="00:02:21.94" heatid="54004" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1156" eventid="30" swimtime="00:01:00.57" lane="1" heatid="30006" points="490">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1157" eventid="34" swimtime="00:01:03.68" lane="2" heatid="34005" points="463">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1158" eventid="42" swimtime="00:00:27.21" lane="2" heatid="42008" points="510" />
                <RESULT resultid="1159" eventid="54" swimtime="00:02:21.47" lane="1" heatid="54004" points="465">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:50.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="265" birthdate="2003-01-01" gender="M" lastname="Reiher" firstname="Janik" license="298654" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:23.56" heatid="44017" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:26.25" heatid="42009" lane="3" />
                <ENTRY eventid="70" entrytime="00:00:23.91" heatid="70001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1160" eventid="44" swimtime="00:00:23.91" lane="1" heatid="44017" points="599" />
                <RESULT resultid="1161" eventid="42" swimtime="00:00:26.20" lane="3" heatid="42009" points="572" />
                <RESULT resultid="2313" eventid="70" swimtime="00:00:23.66" lane="1" heatid="70001" points="618" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="266" birthdate="2015-01-01" gender="F" lastname="Tamm" firstname="Charlotte" license="467460" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.45" heatid="3014" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:38.00" heatid="7019" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:47.31" heatid="13006" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:48.12" heatid="17013" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1162" eventid="3" swimtime="00:00:44.10" lane="2" heatid="3014" points="187" />
                <RESULT resultid="1163" eventid="7" swimtime="00:00:35.71" lane="4" heatid="7019" points="264" />
                <RESULT resultid="1164" eventid="13" swimtime="00:00:47.08" lane="2" heatid="13006" points="138" />
                <RESULT resultid="1165" eventid="17" swimtime="00:00:49.48" lane="4" heatid="17013" points="188" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="KLUB PLAVCÙ MÌLNICKÝCH" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="37" birthdate="2011-01-01" gender="M" lastname="URNER" firstname="DANIEL" license="63439457">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:33.32" heatid="44002" lane="2" />
                <ENTRY eventid="48" entrytime="00:01:22.24" heatid="48003" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:37.76" heatid="26002" lane="2" />
                <ENTRY eventid="32" entrytime="00:01:15.19" heatid="32002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="137" eventid="44" status="DNS" swimtime="00:00:00.00" lane="2" heatid="44002" />
                <RESULT resultid="138" eventid="48" swimtime="00:01:20.33" lane="4" heatid="48003" points="217">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="139" eventid="26" swimtime="00:00:35.92" lane="2" heatid="26002" points="233" />
                <RESULT resultid="177" eventid="32" swimtime="00:01:15.86" lane="1" heatid="32002" points="206">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="39" birthdate="2009-01-01" gender="F" lastname="STRUPLOVÁ" firstname="ELLEN" license="63198000">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:32.71" heatid="43005" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:25.50" heatid="47002" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:38.76" heatid="25002" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:09.18" heatid="31007" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="141" eventid="43" swimtime="00:00:33.97" lane="3" heatid="43005" points="307" />
                <RESULT resultid="142" eventid="47" swimtime="00:01:26.51" lane="3" heatid="47002" points="255">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="143" eventid="25" swimtime="00:00:42.08" lane="2" heatid="25002" points="216" />
                <RESULT resultid="144" eventid="31" swimtime="00:01:12.37" lane="1" heatid="31007" points="334">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="40" birthdate="2010-01-01" gender="M" lastname="MATOUSEK" firstname="JAKUB" license="63461491">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.30" heatid="44010" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:33.75" heatid="28006" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:08.05" heatid="34007" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:29.11" heatid="42005" lane="2" />
                <ENTRY eventid="46" entrytime="00:01:17.61" heatid="46003" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:01.18" heatid="32006" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="145" eventid="44" swimtime="00:00:26.39" lane="4" heatid="44010" points="445" />
                <RESULT resultid="146" eventid="28" swimtime="00:00:33.27" lane="1" heatid="28006" points="421" />
                <RESULT resultid="147" eventid="34" swimtime="00:01:07.42" lane="4" heatid="34007" points="390">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="148" eventid="42" swimtime="00:00:28.84" lane="2" heatid="42005" points="428" />
                <RESULT resultid="149" eventid="46" swimtime="00:01:14.52" lane="4" heatid="46003" points="408">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="150" eventid="32" swimtime="00:00:59.11" lane="3" heatid="32006" points="436">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="41" birthdate="2008-01-01" gender="F" lastname="PETRZELKOVÁ" firstname="JULIE" license="63230000">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:35.19" heatid="43000" lane="0" />
                <ENTRY eventid="25" entrytime="00:00:43.91" heatid="25000" lane="0" />
                <ENTRY eventid="31" entrytime="00:01:19.62" heatid="31000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="151" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
                <RESULT resultid="152" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
                <RESULT resultid="153" eventid="31" status="WDR" swimtime="00:00:00.00" lane="0" heatid="31000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="42" birthdate="2007-01-01" gender="F" lastname="ZLOSKÁ" firstname="KAROLÍNA" license="50882000">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.99" heatid="43013" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:19.01" heatid="33009" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:34.12" heatid="41011" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:08.90" heatid="31012" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="154" eventid="43" swimtime="00:00:31.59" lane="4" heatid="43013" points="382" />
                <RESULT resultid="155" eventid="33" swimtime="00:01:21.53" lane="1" heatid="33009" points="332">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="156" eventid="41" swimtime="00:00:35.25" lane="4" heatid="41011" points="330" />
                <RESULT resultid="157" eventid="31" swimtime="00:01:10.73" lane="1" heatid="31012" points="358">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="43" birthdate="2010-01-01" gender="F" lastname="NOVÁ" firstname="KLÁRA" license="63435167">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:32.31" heatid="43006" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:43.19" heatid="27004" lane="4" />
                <ENTRY eventid="25" entrytime="00:00:38.26" heatid="25003" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:12.55" heatid="31005" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="158" eventid="43" swimtime="00:00:31.25" lane="4" heatid="43006" points="395" />
                <RESULT resultid="159" eventid="27" swimtime="00:00:44.28" lane="4" heatid="27004" points="262" />
                <RESULT resultid="160" eventid="25" swimtime="00:00:39.92" lane="4" heatid="25003" points="253" />
                <RESULT resultid="161" eventid="31" swimtime="00:01:17.91" lane="2" heatid="31005" points="268">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2009-01-01" gender="M" lastname="ZAPP" firstname="MAX" license="63443330">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:26.76" heatid="44000" lane="0" />
                <ENTRY eventid="28" entrytime="00:00:33.45" heatid="28000" lane="0" />
                <ENTRY eventid="38" entrytime="00:02:40.47" heatid="38000" lane="0" />
                <ENTRY eventid="46" entrytime="00:01:13.07" heatid="46000" lane="0" />
                <ENTRY eventid="32" entrytime="00:00:59.12" heatid="32000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="162" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="163" eventid="28" status="WDR" swimtime="00:00:00.00" lane="0" heatid="28000" />
                <RESULT resultid="164" eventid="38" status="WDR" swimtime="00:00:00.00" lane="0" heatid="38000" />
                <RESULT resultid="165" eventid="46" status="WDR" swimtime="00:00:00.00" lane="0" heatid="46000" />
                <RESULT resultid="166" eventid="32" status="WDR" swimtime="00:00:00.00" lane="0" heatid="32000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="45" birthdate="2011-01-01" gender="F" lastname="TESÁRKOVÁ" firstname="PAVLÍNA" license="63455188">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:35.17" heatid="43003" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:43.59" heatid="27003" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:32.78" heatid="33002" lane="1" />
                <ENTRY eventid="45" entrytime="00:01:33.75" heatid="45005" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:19.75" heatid="31002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="167" eventid="43" swimtime="00:00:34.58" lane="1" heatid="43003" points="291" />
                <RESULT resultid="168" eventid="27" swimtime="00:00:42.55" lane="3" heatid="27003" points="296" />
                <RESULT resultid="169" eventid="33" swimtime="00:01:28.22" lane="1" heatid="33002" points="262">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="170" eventid="45" swimtime="00:01:33.56" lane="4" heatid="45005" points="296">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="171" eventid="31" swimtime="00:01:18.03" lane="2" heatid="31002" points="267">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="46" birthdate="2010-01-01" gender="M" lastname="ZNAMENÁÈEK" firstname="STÌPÁN" license="63465074">
              <ENTRIES>
                <ENTRY eventid="32" entrytime="00:01:12.58" heatid="32002" lane="2" />
                <ENTRY eventid="44" entrytime="00:00:32.04" heatid="44003" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:41.25" heatid="28003" lane="4" />
                <ENTRY eventid="34" entrytime="00:01:26.41" heatid="34001" lane="3" />
                <ENTRY eventid="46" entrytime="00:01:28.95" heatid="46001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="172" eventid="44" status="DNS" swimtime="00:00:00.00" lane="3" heatid="44003" />
                <RESULT resultid="173" eventid="28" status="DSQ" swimtime="00:00:41.13" lane="4" heatid="28003" comment="Nach dem Start hat der Sportler zwei Delphinbeinschläge ausgeführt." />
                <RESULT resultid="174" eventid="34" swimtime="00:01:22.64" lane="3" heatid="34001" points="212">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="175" eventid="46" swimtime="00:01:28.15" lane="3" heatid="46001" points="246">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="176" eventid="32" swimtime="00:01:12.91" lane="2" heatid="32002" points="232">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="KS Swim Team Nowa Ruda" nation="POL" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="267" birthdate="2011-01-01" gender="F" lastname="Cergier" firstname="Samanta" license="0">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:35.40" heatid="43002" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:44.20" heatid="27003" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:21.10" heatid="33007" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1166" eventid="43" swimtime="00:00:37.09" lane="2" heatid="43002" points="236" />
                <RESULT resultid="1167" eventid="27" swimtime="00:00:47.68" lane="4" heatid="27003" points="210" />
                <RESULT resultid="1168" eventid="33" status="DSQ" swimtime="00:01:32.66" lane="1" heatid="33007" comment="Die Teilstrecke Rücken wurde nicht in Rückenlage beendet.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="268" birthdate="2013-01-01" gender="F" lastname="Mostowy" firstname="Maja" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:46.10" heatid="3013" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:22.10" heatid="19018" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1169" eventid="3" swimtime="00:00:41.43" lane="2" heatid="3013" points="226" />
                <RESULT resultid="1170" eventid="19" swimtime="00:01:27.18" lane="1" heatid="19018" points="191">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="269" birthdate="2017-01-01" gender="F" lastname="Mostowy" firstname="Martyna" license="0">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:00:51.00" heatid="7006" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:57.10" heatid="17016" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1171" eventid="7" swimtime="00:00:48.24" lane="4" heatid="7006" points="107" />
                <RESULT resultid="1172" eventid="17" swimtime="00:01:02.19" lane="4" heatid="17016" points="94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="270" birthdate="2016-01-01" gender="F" lastname="Pasek" firstname="Laura" license="0">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:45.00" heatid="5012" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:41.00" heatid="7014" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:48.10" heatid="17017" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1173" eventid="5" swimtime="00:01:52.90" lane="3" heatid="5012" points="168">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1174" eventid="7" swimtime="00:00:41.93" lane="2" heatid="7014" points="163" />
                <RESULT resultid="1175" eventid="17" swimtime="00:00:48.89" lane="3" heatid="17017" points="195" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="271" birthdate="2011-01-01" gender="F" lastname="Ryskiewicz" firstname="Maja" license="0">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:37.80" heatid="43001" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:31.80" heatid="47001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1176" eventid="43" swimtime="00:00:43.03" lane="3" heatid="43001" points="151" />
                <RESULT resultid="1177" eventid="47" swimtime="00:01:48.12" lane="2" heatid="47001" points="130">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Neratovicky plavecky klub" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="153" birthdate="2015-01-01" gender="M" lastname="Cerny" firstname="Radek" license="0">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:42.39" heatid="2003" lane="3" />
                <ENTRY eventid="6" entrytime="00:01:36.65" heatid="6009" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:34.62" heatid="8022" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:43.94" heatid="18012" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:19.16" heatid="20019" lane="1" />
                <ENTRY eventid="22" entrytime="00:03:10.90" heatid="22000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="705" eventid="2" status="DNS" swimtime="00:00:00.00" lane="3" heatid="2003" />
                <RESULT resultid="706" eventid="6" status="DNS" swimtime="00:00:00.00" lane="4" heatid="6009" />
                <RESULT resultid="707" eventid="8" status="WDR" swimtime="00:00:00.00" lane="1" heatid="8022" />
                <RESULT resultid="708" eventid="18" status="WDR" swimtime="00:00:00.00" lane="1" heatid="18012" />
                <RESULT resultid="709" eventid="20" status="WDR" swimtime="00:00:00.00" lane="1" heatid="20019" />
                <RESULT resultid="710" eventid="22" status="WDR" swimtime="00:00:00.00" lane="0" heatid="22000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154" birthdate="2015-01-01" gender="F" lastname="Filipkova" firstname="Kristyna" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:52.26" heatid="3008" lane="2" />
                <ENTRY eventid="5" entrytime="00:01:50.21" heatid="5006" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:44.01" heatid="7011" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:51.01" heatid="17010" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:43.17" heatid="19008" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="711" eventid="3" status="DNS" swimtime="00:00:00.00" lane="2" heatid="3008" />
                <RESULT resultid="712" eventid="5" status="DNS" swimtime="00:00:00.00" lane="1" heatid="5006" />
                <RESULT resultid="713" eventid="7" status="DNS" swimtime="00:00:00.00" lane="2" heatid="7011" />
                <RESULT resultid="714" eventid="17" status="DNS" swimtime="00:00:00.00" lane="3" heatid="17010" />
                <RESULT resultid="715" eventid="19" status="DNS" swimtime="00:00:00.00" lane="1" heatid="19008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="155" birthdate="2015-01-01" gender="F" lastname="Franova" firstname="Zita" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.00" heatid="3015" lane="3" />
                <ENTRY eventid="5" entrytime="00:01:47.69" heatid="5007" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:35.82" heatid="7023" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:40.23" heatid="15009" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:48.16" heatid="17012" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:22.32" heatid="19018" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="716" eventid="3" swimtime="00:00:44.21" lane="3" heatid="3015" points="186" />
                <RESULT resultid="717" eventid="5" swimtime="00:01:49.75" lane="4" heatid="5007" points="183">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="718" eventid="7" swimtime="00:00:35.83" lane="1" heatid="7023" points="262" />
                <RESULT resultid="719" eventid="15" swimtime="00:01:37.11" lane="1" heatid="15009" points="180">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="720" eventid="17" swimtime="00:00:50.04" lane="2" heatid="17012" points="182" />
                <RESULT resultid="721" eventid="19" swimtime="00:01:19.53" lane="4" heatid="19018" points="252">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156" birthdate="2012-01-01" gender="M" lastname="Kouba" firstname="Daniel" license="0">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:46.83" heatid="2001" lane="3" />
                <ENTRY eventid="6" entrytime="00:01:39.47" heatid="6006" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:36.41" heatid="8013" lane="1" />
                <ENTRY eventid="16" entrytime="00:01:39.80" heatid="16004" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:46.48" heatid="18007" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:19.86" heatid="20012" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="722" eventid="2" swimtime="00:01:40.45" lane="3" heatid="2001" points="107">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="723" eventid="6" swimtime="00:01:43.70" lane="1" heatid="6006" points="151">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="724" eventid="8" swimtime="00:00:35.62" lane="1" heatid="8013" points="181" />
                <RESULT resultid="725" eventid="16" swimtime="00:01:45.67" lane="1" heatid="16004" points="95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="726" eventid="18" swimtime="00:00:46.97" lane="3" heatid="18007" points="149" />
                <RESULT resultid="727" eventid="20" swimtime="00:01:18.64" lane="3" heatid="20012" points="185">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157" birthdate="2013-01-01" gender="F" lastname="Poddana" firstname="Viktorie" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:42.09" heatid="3017" lane="3" />
                <ENTRY eventid="5" entrytime="00:01:45.52" heatid="5007" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:34.99" heatid="7024" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:36.11" heatid="15011" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:49.54" heatid="17011" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:19.57" heatid="19020" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="728" eventid="3" swimtime="00:00:39.63" lane="3" heatid="3017" points="258" />
                <RESULT resultid="729" eventid="5" swimtime="00:01:46.64" lane="2" heatid="5007" points="199">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="730" eventid="7" swimtime="00:00:33.81" lane="4" heatid="7024" points="311" />
                <RESULT resultid="731" eventid="15" swimtime="00:01:29.42" lane="1" heatid="15011" points="231">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="732" eventid="17" swimtime="00:00:50.20" lane="3" heatid="17011" points="180" />
                <RESULT resultid="733" eventid="19" swimtime="00:01:16.89" lane="4" heatid="19020" points="279">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="158" birthdate="2016-01-01" gender="M" lastname="Schurmann" firstname="Oliver" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:58.42" heatid="4002" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:50.37" heatid="8003" lane="2" />
                <ENTRY eventid="18" entrytime="00:01:00.27" heatid="18002" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:54.65" heatid="20002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="734" eventid="4" swimtime="00:00:55.30" lane="4" heatid="4002" points="63" />
                <RESULT resultid="735" eventid="8" swimtime="00:00:44.61" lane="2" heatid="8003" points="92" />
                <RESULT resultid="736" eventid="18" swimtime="00:00:57.88" lane="2" heatid="18002" points="80" />
                <RESULT resultid="737" eventid="20" swimtime="00:01:45.21" lane="2" heatid="20002" points="77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="159" birthdate="2016-01-01" gender="F" lastname="Skruzna" firstname="Laura" license="0">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:58.76" heatid="5000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:48.90" heatid="7000" lane="0" />
                <ENTRY eventid="17" entrytime="00:00:52.35" heatid="17000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:50.60" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="738" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="739" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="740" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
                <RESULT resultid="741" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2016-01-01" gender="M" lastname="Skruzny" firstname="Daniel" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:51.47" heatid="6000" lane="0" />
                <ENTRY eventid="8" entrytime="00:00:43.77" heatid="8000" lane="0" />
                <ENTRY eventid="18" entrytime="00:00:51.53" heatid="18000" lane="0" />
                <ENTRY eventid="20" entrytime="00:01:42.45" heatid="20000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="742" eventid="6" status="WDR" swimtime="00:00:00.00" lane="0" heatid="6000" />
                <RESULT resultid="743" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="744" eventid="18" status="WDR" swimtime="00:00:00.00" lane="0" heatid="18000" />
                <RESULT resultid="745" eventid="20" status="WDR" swimtime="00:00:00.00" lane="0" heatid="20000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2013-01-01" gender="M" lastname="Tomasek" firstname="Dan" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:26.45" heatid="6000" lane="0" />
                <ENTRY eventid="8" entrytime="00:00:31.19" heatid="8000" lane="0" />
                <ENTRY eventid="10" entrytime="00:01:19.24" heatid="10000" lane="0" />
                <ENTRY eventid="18" entrytime="00:00:38.17" heatid="18000" lane="0" />
                <ENTRY eventid="20" entrytime="00:01:11.25" heatid="20000" lane="0" />
                <ENTRY eventid="22" entrytime="00:02:54.12" heatid="22000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="746" eventid="6" status="WDR" swimtime="00:00:00.00" lane="0" heatid="6000" />
                <RESULT resultid="747" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="748" eventid="10" status="WDR" swimtime="00:00:00.00" lane="0" heatid="10000" />
                <RESULT resultid="749" eventid="18" status="WDR" swimtime="00:00:00.00" lane="0" heatid="18000" />
                <RESULT resultid="750" eventid="20" status="WDR" swimtime="00:00:00.00" lane="0" heatid="20000" />
                <RESULT resultid="751" eventid="22" status="WDR" swimtime="00:00:00.00" lane="0" heatid="22000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="162" birthdate="2016-01-01" gender="M" lastname="Tvrdik" firstname="Daniel" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:02:04.22" heatid="6002" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:56.26" heatid="8001" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:57.98" heatid="18003" lane="1" />
                <ENTRY eventid="20" entrytime="00:02:02.06" heatid="20002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="752" eventid="6" swimtime="00:02:10.30" lane="1" heatid="6002" points="76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="753" eventid="8" swimtime="00:00:51.73" lane="2" heatid="8001" points="59" />
                <RESULT resultid="754" eventid="18" swimtime="00:00:59.24" lane="1" heatid="18003" points="74" />
                <RESULT resultid="755" eventid="20" swimtime="00:01:54.33" lane="4" heatid="20002" points="60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163" birthdate="2014-01-01" gender="M" lastname="Tvrdik" firstname="Matteo" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:44.29" heatid="6010" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:34.26" heatid="8016" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:34.09" heatid="10004" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:48.30" heatid="18013" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:18.75" heatid="20012" lane="2" />
                <ENTRY eventid="22" entrytime="00:03:23.49" heatid="22002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="756" eventid="6" status="DNS" swimtime="00:00:00.00" lane="1" heatid="6010" />
                <RESULT resultid="757" eventid="8" status="DNS" swimtime="00:00:00.00" lane="2" heatid="8016" />
                <RESULT resultid="758" eventid="10" status="DNS" swimtime="00:00:00.00" lane="2" heatid="10004" />
                <RESULT resultid="759" eventid="18" status="DNS" swimtime="00:00:00.00" lane="4" heatid="18013" />
                <RESULT resultid="760" eventid="20" status="DNS" swimtime="00:00:00.00" lane="2" heatid="20012" />
                <RESULT resultid="761" eventid="22" status="DNS" swimtime="00:00:00.00" lane="3" heatid="22002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Plavecký klub Litvínov" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="119" birthdate="2016-01-01" gender="F" lastname="HAASOVÁ" firstname="Veronika" license="63454639">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:02:03.65" heatid="5003" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:41.86" heatid="7014" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:48.86" heatid="13005" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:54.34" heatid="17007" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="562" eventid="5" swimtime="00:02:04.52" lane="3" heatid="5003" points="125">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="563" eventid="7" swimtime="00:00:42.74" lane="4" heatid="7014" points="154" />
                <RESULT resultid="564" eventid="13" swimtime="00:00:47.04" lane="4" heatid="13005" points="139" />
                <RESULT resultid="565" eventid="17" swimtime="00:00:56.17" lane="3" heatid="17007" points="128" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120" birthdate="2016-01-01" gender="M" lastname="JANDOVSKÝ" firstname="Stepán" license="63459278">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:00:35.68" heatid="8021" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:33.06" heatid="10009" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:42.47" heatid="14008" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:42.21" heatid="16007" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="566" eventid="8" swimtime="00:00:36.07" lane="2" heatid="8021" points="174" />
                <RESULT resultid="567" eventid="10" swimtime="00:01:31.50" lane="2" heatid="10009" points="156">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="568" eventid="14" swimtime="00:00:42.96" lane="2" heatid="14008" points="129" />
                <RESULT resultid="569" eventid="16" swimtime="00:01:31.90" lane="4" heatid="16007" points="145">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121" birthdate="2016-01-01" gender="M" lastname="KOMLÓ" firstname="Jakub Michal" license="63459269">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:45.27" heatid="4000" lane="0" />
                <ENTRY eventid="6" entrytime="00:01:49.19" heatid="6000" lane="0" />
                <ENTRY eventid="18" entrytime="00:00:50.55" heatid="18000" lane="0" />
                <ENTRY eventid="20" entrytime="00:01:36.17" heatid="20000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="570" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="571" eventid="6" status="WDR" swimtime="00:00:00.00" lane="0" heatid="6000" />
                <RESULT resultid="572" eventid="18" status="WDR" swimtime="00:00:00.00" lane="0" heatid="18000" />
                <RESULT resultid="573" eventid="20" status="WDR" swimtime="00:00:00.00" lane="0" heatid="20000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122" birthdate="2017-01-01" gender="M" lastname="KORÍNEK" firstname="Tomás" license="63454638">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:50.12" heatid="4000" lane="0" />
                <ENTRY eventid="8" entrytime="00:00:43.61" heatid="8000" lane="0" />
                <ENTRY eventid="16" entrytime="00:01:47.40" heatid="16000" lane="0" />
                <ENTRY eventid="20" entrytime="00:01:43.09" heatid="20000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="574" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="575" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="576" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="577" eventid="20" status="WDR" swimtime="00:00:00.00" lane="0" heatid="20000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123" birthdate="2014-01-01" gender="F" lastname="KUKANOVÁ" firstname="Sára" license="63474909">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:46.82" heatid="3000" lane="0" />
                <ENTRY eventid="9" entrytime="00:01:44.43" heatid="9000" lane="0" />
                <ENTRY eventid="15" entrytime="00:01:38.76" heatid="15000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:27.44" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="578" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="579" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
                <RESULT resultid="580" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="581" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124" birthdate="2013-01-01" gender="F" lastname="LANGHAMMEROVÁ" firstname="Ella" license="63459214">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:42.29" heatid="5009" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:36.14" heatid="7022" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:47.13" heatid="17013" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:21.08" heatid="19019" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="582" eventid="5" status="DNS" swimtime="00:00:00.00" lane="2" heatid="5009" />
                <RESULT resultid="583" eventid="7" status="DNS" swimtime="00:00:00.00" lane="2" heatid="7022" />
                <RESULT resultid="584" eventid="17" status="DNS" swimtime="00:00:00.00" lane="2" heatid="17013" />
                <RESULT resultid="585" eventid="19" status="DNS" swimtime="00:00:00.00" lane="3" heatid="19019" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125" birthdate="2016-01-01" gender="M" lastname="LENCÉS" firstname="Jan" license="63467350">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:48.63" heatid="4007" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:41.60" heatid="8009" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:57.12" heatid="18003" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:39.23" heatid="20005" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="586" eventid="4" swimtime="00:00:46.59" lane="4" heatid="4007" points="106" />
                <RESULT resultid="587" eventid="8" swimtime="00:00:40.50" lane="4" heatid="8009" points="123" />
                <RESULT resultid="588" eventid="18" swimtime="00:00:58.64" lane="2" heatid="18003" points="77" />
                <RESULT resultid="589" eventid="20" swimtime="00:01:36.72" lane="4" heatid="20005" points="99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="126" birthdate="2016-01-01" gender="F" lastname="ULRICHOVÁ" firstname="Anezka" license="63454648">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:47.30" heatid="3012" lane="1" />
                <ENTRY eventid="5" entrytime="00:01:41.41" heatid="5012" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:42.90" heatid="15016" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:34.54" heatid="19011" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="590" eventid="3" swimtime="00:00:45.60" lane="1" heatid="3012" points="169" />
                <RESULT resultid="591" eventid="5" swimtime="00:01:56.57" lane="2" heatid="5012" points="153">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="592" eventid="15" swimtime="00:01:40.31" lane="4" heatid="15016" points="163">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="593" eventid="19" swimtime="00:01:32.46" lane="3" heatid="19011" points="160">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="127" birthdate="2015-01-01" gender="F" lastname="VOJTULOVICOVÁ" firstname="Ema" license="63454640">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:46.42" heatid="3013" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:37.90" heatid="7019" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:45.60" heatid="13007" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:39.14" heatid="15010" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="594" eventid="3" status="DSQ" swimtime="00:00:45.77" lane="1" heatid="3013" comment="Die Sportlerin hat bei der Wende nach Verlassen der Rückenlage nicht unverzüglich die eigentliche Wendenbewegung ausgeführt." />
                <RESULT resultid="595" eventid="7" swimtime="00:00:38.16" lane="1" heatid="7019" points="216" />
                <RESULT resultid="596" eventid="13" swimtime="00:00:44.68" lane="3" heatid="13007" points="162" />
                <RESULT resultid="597" eventid="15" swimtime="00:01:40.67" lane="4" heatid="15010" points="162">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:01:51.81" lane="0" heatid="11000" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="561" eventid="11" status="WDR" swimtime="00:00:00.00" lane="0" heatid="11000" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Plavecký klub Most" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="104" birthdate="2010-01-01" gender="M" lastname="Augustín" firstname="Tomas" license="0">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:26.99" heatid="44010" lane="2" />
                <ENTRY eventid="34" entrytime="00:01:08.48" heatid="34005" lane="1" />
                <ENTRY eventid="52" entrytime="00:02:10.78" heatid="52004" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:28.55" heatid="42007" lane="3" />
                <ENTRY eventid="32" entrytime="00:00:58.76" heatid="32011" lane="4" />
                <ENTRY eventid="54" entrytime="00:02:28.92" heatid="54003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="493" eventid="44" swimtime="00:00:26.82" lane="2" heatid="44010" points="424" />
                <RESULT resultid="494" eventid="34" swimtime="00:01:10.25" lane="1" heatid="34005" points="345">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="495" eventid="52" swimtime="00:02:17.14" lane="2" heatid="52004" points="380">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:06.87" />
                    <SPLIT distance="150" swimtime="00:01:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="496" eventid="42" swimtime="00:00:29.35" lane="3" heatid="42007" points="406" />
                <RESULT resultid="497" eventid="32" swimtime="00:01:02.71" lane="4" heatid="32011" points="365">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="498" eventid="54" swimtime="00:02:40.18" lane="1" heatid="54003" points="320">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="150" swimtime="00:01:59.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105" birthdate="2016-01-01" gender="F" lastname="Berkyová" firstname="Victoria" license="0">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:00:38.10" heatid="7018" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:47.10" heatid="9004" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:48.00" heatid="13006" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:26.98" heatid="19022" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="499" eventid="7" swimtime="00:00:37.71" lane="3" heatid="7018" points="224" />
                <RESULT resultid="500" eventid="9" swimtime="00:01:44.01" lane="1" heatid="9004" points="160">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="501" eventid="13" swimtime="00:00:51.64" lane="4" heatid="13006" points="105" />
                <RESULT resultid="502" eventid="19" swimtime="00:01:26.18" lane="4" heatid="19022" points="198">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106" birthdate="2014-01-01" gender="F" lastname="Bulei" firstname="Daryna" license="0">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:50.62" heatid="1001" lane="1" />
                <ENTRY eventid="5" entrytime="00:01:49.77" heatid="5006" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:36.77" heatid="9008" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:36.30" heatid="15011" lane="4" />
                <ENTRY eventid="21" entrytime="00:03:23.78" heatid="21001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="503" eventid="1" swimtime="00:01:47.82" lane="1" heatid="1001" points="125">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="504" eventid="5" swimtime="00:01:46.78" lane="3" heatid="5006" points="199">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="505" eventid="9" swimtime="00:01:34.15" lane="1" heatid="9008" points="216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="506" eventid="15" swimtime="00:01:34.56" lane="4" heatid="15011" points="195">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="507" eventid="21" swimtime="00:03:22.13" lane="2" heatid="21001" points="219">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                    <SPLIT distance="100" swimtime="00:01:38.73" />
                    <SPLIT distance="150" swimtime="00:02:36.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="2013-01-01" gender="M" lastname="Capek" firstname="Tomás" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:42.94" heatid="4009" lane="3" />
                <ENTRY eventid="6" entrytime="00:01:45.61" heatid="6005" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:36.03" heatid="8013" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:33.26" heatid="16010" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:16.68" heatid="20013" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="508" eventid="4" swimtime="00:00:44.55" lane="3" heatid="4009" points="122" />
                <RESULT resultid="509" eventid="6" swimtime="00:01:46.36" lane="1" heatid="6005" points="140">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="510" eventid="8" swimtime="00:00:36.92" lane="2" heatid="8013" points="162" />
                <RESULT resultid="511" eventid="16" status="DSQ" swimtime="00:01:33.03" lane="4" heatid="16010" comment="Bei der zweiten Wende hat der Sportler die Wand verlassen, bevor die Rückenlage eingenommen war.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="512" eventid="20" swimtime="00:01:17.97" lane="3" heatid="20013" points="190">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2010-01-01" gender="M" lastname="Fedori" firstname="Daniil" license="0">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.66" heatid="44007" lane="2" />
                <ENTRY eventid="30" entrytime="00:01:10.14" heatid="30002" lane="1" />
                <ENTRY eventid="48" entrytime="00:01:06.83" heatid="48004" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:29.01" heatid="42006" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:30.63" heatid="26008" lane="1" />
                <ENTRY eventid="36" entrytime="00:02:31.11" heatid="36002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="513" eventid="44" swimtime="00:00:27.82" lane="2" heatid="44007" points="380" />
                <RESULT resultid="514" eventid="30" swimtime="00:01:08.17" lane="1" heatid="30002" points="344">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="515" eventid="48" swimtime="00:01:07.98" lane="1" heatid="48004" points="359">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="516" eventid="42" swimtime="00:00:28.80" lane="3" heatid="42006" points="430" />
                <RESULT resultid="517" eventid="26" swimtime="00:00:30.03" lane="1" heatid="26008" points="399" />
                <RESULT resultid="518" eventid="36" swimtime="00:02:27.98" lane="1" heatid="36002" points="363">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="150" swimtime="00:01:53.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="2013-01-01" gender="F" lastname="Kolariková" firstname="Nikola" license="0">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:45.00" heatid="5008" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:35.70" heatid="9009" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:47.71" heatid="13006" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:26.14" heatid="19015" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="519" eventid="5" swimtime="00:01:43.92" lane="1" heatid="5008" points="216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="520" eventid="9" swimtime="00:01:34.50" lane="1" heatid="9009" points="213">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="521" eventid="13" swimtime="00:00:46.28" lane="1" heatid="13006" points="146" />
                <RESULT resultid="522" eventid="19" swimtime="00:01:26.31" lane="4" heatid="19015" points="197">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110" birthdate="2010-01-01" gender="F" lastname="Komínková" firstname="Pavlína" license="0">
              <ENTRIES>
                <ENTRY eventid="37" entrytime="00:02:39.88" heatid="37002" lane="3" />
                <ENTRY eventid="53" entrytime="00:02:29.63" heatid="53003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="523" eventid="37" swimtime="00:02:41.92" lane="3" heatid="37002" points="574">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:18.48" />
                    <SPLIT distance="150" swimtime="00:02:00.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="524" eventid="53" swimtime="00:02:30.00" lane="3" heatid="53003" points="536">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:52.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111" birthdate="2017-01-01" gender="M" lastname="Kuranda" firstname="Tobias" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:53.84" heatid="4011" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:45.34" heatid="8020" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:58.19" heatid="16006" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:43.49" heatid="20017" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="525" eventid="4" swimtime="00:00:51.78" lane="2" heatid="4011" points="77" />
                <RESULT resultid="526" eventid="8" swimtime="00:00:45.05" lane="3" heatid="8020" points="89" />
                <RESULT resultid="527" eventid="16" status="DSQ" swimtime="00:01:51.84" lane="4" heatid="16006" comment="Der Sportler hat bei der ersten Wende nach Verlassen der Rückenlage nicht unverzüglich die eigentliche Wendenbewegung ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="528" eventid="20" swimtime="00:01:39.95" lane="3" heatid="20017" points="90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="112" birthdate="2015-01-01" gender="M" lastname="Martínek" firstname="Jan" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:36.63" heatid="6009" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:34.61" heatid="8022" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:25.85" heatid="10010" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:42.51" heatid="14009" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:16.57" heatid="20019" lane="2" />
                <ENTRY eventid="22" entrytime="00:03:17.11" heatid="22003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="529" eventid="6" swimtime="00:01:35.84" lane="1" heatid="6009" points="191">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="530" eventid="8" swimtime="00:00:35.19" lane="3" heatid="8022" points="188" />
                <RESULT resultid="531" eventid="10" swimtime="00:01:26.49" lane="2" heatid="10010" points="184">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="532" eventid="14" swimtime="00:00:45.28" lane="2" heatid="14009" points="110" />
                <RESULT resultid="533" eventid="20" swimtime="00:01:15.89" lane="2" heatid="20019" points="206">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="534" eventid="22" swimtime="00:03:10.79" lane="4" heatid="22003" points="189">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.45" />
                    <SPLIT distance="100" swimtime="00:01:35.59" />
                    <SPLIT distance="150" swimtime="00:02:28.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113" birthdate="2009-01-01" gender="M" lastname="Najmon" firstname="Tomás" license="0">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:33.89" heatid="28006" lane="4" />
                <ENTRY eventid="34" entrytime="00:01:07.54" heatid="34007" lane="1" />
                <ENTRY eventid="38" entrytime="00:02:47.51" heatid="38005" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:12.93" heatid="46005" lane="4" />
                <ENTRY eventid="54" entrytime="00:02:25.39" heatid="54003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="535" eventid="28" swimtime="00:00:34.20" lane="4" heatid="28006" points="388" />
                <RESULT resultid="536" eventid="34" swimtime="00:01:09.07" lane="1" heatid="34007" points="363">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="537" eventid="38" swimtime="00:02:49.66" lane="4" heatid="38005" points="355">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:06.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="538" eventid="46" swimtime="00:01:15.26" lane="4" heatid="46005" points="396">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="539" eventid="54" swimtime="00:02:27.43" lane="2" heatid="54003" points="411">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:11.72" />
                    <SPLIT distance="150" swimtime="00:01:53.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="114" birthdate="2012-01-01" gender="F" lastname="Rejmanová" firstname="Laura" license="0">
              <ENTRIES>
                <ENTRY eventid="47" entrytime="00:01:55.09" heatid="47001" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:55.00" heatid="33001" lane="1" />
                <ENTRY eventid="25" entrytime="00:00:54.44" heatid="25001" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:44.07" heatid="31001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="540" eventid="47" swimtime="00:01:49.86" lane="4" heatid="47001" points="124">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="541" eventid="33" swimtime="00:01:52.69" lane="1" heatid="33001" points="126">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="542" eventid="25" swimtime="00:00:49.16" lane="4" heatid="25001" points="135" />
                <RESULT resultid="543" eventid="31" status="DSQ" swimtime="00:01:41.60" lane="1" heatid="31001" comment="Bei der dritten Wende wurde die Wand nicht berührt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="115" birthdate="2014-01-01" gender="M" lastname="Rychly" firstname="Jan" license="0">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:14.33" heatid="2004" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:29.75" heatid="8023" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:13.27" heatid="10011" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:31.93" heatid="14010" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:05.01" heatid="20020" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="544" eventid="2" swimtime="00:01:15.40" lane="2" heatid="2004" points="254">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="545" eventid="8" swimtime="00:00:29.12" lane="2" heatid="8023" points="331" />
                <RESULT resultid="546" eventid="10" swimtime="00:01:14.11" lane="2" heatid="10011" points="294">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="547" eventid="14" swimtime="00:00:31.78" lane="2" heatid="14010" points="320" />
                <RESULT resultid="548" eventid="20" swimtime="00:01:05.44" lane="2" heatid="20020" points="321">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="116" birthdate="2014-01-01" gender="M" lastname="Vacek" firstname="Jachym" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:37.80" heatid="4014" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:32.32" heatid="8023" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:21.09" heatid="10011" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:35.36" heatid="14010" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:10.20" heatid="20020" lane="3" />
                <ENTRY eventid="22" entrytime="00:02:52.41" heatid="22004" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="549" eventid="4" swimtime="00:00:37.34" lane="3" heatid="4014" points="207" />
                <RESULT resultid="550" eventid="8" swimtime="00:00:31.87" lane="4" heatid="8023" points="253" />
                <RESULT resultid="551" eventid="10" swimtime="00:01:20.89" lane="3" heatid="10011" points="226">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="552" eventid="14" swimtime="00:00:35.88" lane="3" heatid="14010" points="222" />
                <RESULT resultid="553" eventid="20" swimtime="00:01:11.41" lane="3" heatid="20020" points="247">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="554" eventid="22" swimtime="00:02:50.19" lane="2" heatid="22004" points="267">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:01:21.84" />
                    <SPLIT distance="150" swimtime="00:02:12.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="117" birthdate="2014-01-01" gender="M" lastname="Valenta" firstname="Krystof" license="0">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:25.85" heatid="2004" lane="1" />
                <ENTRY eventid="4" entrytime="00:00:38.95" heatid="4014" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:21.71" heatid="10011" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:37.42" heatid="14007" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:19.81" heatid="16009" lane="3" />
                <ENTRY eventid="22" entrytime="00:02:52.44" heatid="22004" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="555" eventid="2" swimtime="00:01:32.08" lane="1" heatid="2004" points="139">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="556" eventid="4" swimtime="00:00:39.65" lane="1" heatid="4014" points="173" />
                <RESULT resultid="557" eventid="10" swimtime="00:01:27.00" lane="1" heatid="10011" points="181">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="558" eventid="14" swimtime="00:00:37.73" lane="3" heatid="14007" points="191" />
                <RESULT resultid="559" eventid="16" swimtime="00:01:22.26" lane="3" heatid="16009" points="202">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="560" eventid="22" swimtime="00:03:03.11" lane="3" heatid="22004" points="214">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                    <SPLIT distance="100" swimtime="00:01:28.53" />
                    <SPLIT distance="150" swimtime="00:02:23.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Chemnitz von 1892" nation="GER" region="12" code="3353">
          <ATHLETES>
            <ATHLETE athleteid="166" birthdate="2011-01-01" gender="M" lastname="Berger" firstname="Paul Alexander" license="448319" nation="GER">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:37.99" heatid="28008" lane="1" />
                <ENTRY eventid="38" entrytime="00:03:02.22" heatid="38004" lane="1" />
                <ENTRY eventid="46" entrytime="00:01:23.37" heatid="46004" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="766" eventid="28" swimtime="00:00:37.47" lane="1" heatid="28008" points="295" />
                <RESULT resultid="767" eventid="38" swimtime="00:03:00.38" lane="1" heatid="38004" points="295">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                    <SPLIT distance="100" swimtime="00:01:28.05" />
                    <SPLIT distance="150" swimtime="00:02:14.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="768" eventid="46" swimtime="00:01:23.76" lane="2" heatid="46004" points="287">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="2011-01-01" gender="F" lastname="Böhm" firstname="Laura" license="423442">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.46" heatid="43011" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:16.12" heatid="33007" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:32.56" heatid="41009" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:08.65" heatid="31010" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="769" eventid="43" swimtime="00:00:29.94" lane="2" heatid="43011" points="449" />
                <RESULT resultid="770" eventid="33" swimtime="00:01:17.04" lane="2" heatid="33007" points="394">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="771" eventid="41" swimtime="00:00:33.42" lane="2" heatid="41009" points="388" />
                <RESULT resultid="772" eventid="31" swimtime="00:01:07.90" lane="3" heatid="31010" points="405">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="168" birthdate="2009-01-01" gender="M" lastname="Degelmann" firstname="Max" license="408969">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:28.15" heatid="44007" lane="1" />
                <ENTRY eventid="48" entrytime="00:01:09.30" heatid="48004" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:31.20" heatid="26008" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:03.30" heatid="32005" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="773" eventid="44" swimtime="00:00:27.77" lane="1" heatid="44007" points="382" />
                <RESULT resultid="774" eventid="48" swimtime="00:01:09.11" lane="4" heatid="48004" points="342">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="775" eventid="26" swimtime="00:00:30.46" lane="4" heatid="26008" points="382" />
                <RESULT resultid="776" eventid="32" swimtime="00:01:02.46" lane="1" heatid="32005" points="369">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169" birthdate="2008-01-01" gender="M" lastname="Gensler" firstname="Daniel" license="365320">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:26.03" heatid="44011" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:32.55" heatid="28010" lane="3" />
                <ENTRY eventid="32" entrytime="00:00:59.08" heatid="32008" lane="2" />
                <ENTRY eventid="61" entrytime="00:00:32.16" heatid="61001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="777" eventid="44" swimtime="00:00:25.44" lane="2" heatid="44011" points="497" />
                <RESULT resultid="778" eventid="28" swimtime="00:00:32.16" lane="3" heatid="28010" points="466" />
                <RESULT resultid="779" eventid="32" swimtime="00:00:56.88" lane="2" heatid="32008" points="489">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2325" eventid="61" swimtime="00:00:31.36" lane="1" heatid="61001" points="503" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170" birthdate="2010-01-01" gender="F" lastname="Gerlach" firstname="Mona" license="413351" nation="GER">
              <ENTRIES>
                <ENTRY eventid="47" entrytime="00:01:17.65" heatid="47003" lane="4" />
                <ENTRY eventid="51" entrytime="00:02:43.27" heatid="51001" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:35.50" heatid="25004" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:10.19" heatid="31006" lane="3" />
                <ENTRY eventid="55" entrytime="00:00:34.75" heatid="55001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="780" eventid="47" swimtime="00:01:15.17" lane="4" heatid="47003" points="389">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="781" eventid="51" swimtime="00:02:29.50" lane="3" heatid="51001" points="401">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:51.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="782" eventid="25" swimtime="00:00:34.75" lane="4" heatid="25004" points="383" />
                <RESULT resultid="783" eventid="31" swimtime="00:01:07.32" lane="3" heatid="31006" points="415">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2350" eventid="55" swimtime="00:00:34.31" lane="4" heatid="55001" points="398" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="171" birthdate="2010-01-01" gender="M" lastname="Hoheisel" firstname="Lukas" license="408976">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.77" heatid="44007" lane="3" />
                <ENTRY eventid="52" entrytime="00:02:30.67" heatid="52003" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:30.57" heatid="42004" lane="2" />
                <ENTRY eventid="32" entrytime="00:01:00.72" heatid="32007" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="784" eventid="44" swimtime="00:00:27.42" lane="3" heatid="44007" points="397" />
                <RESULT resultid="785" eventid="52" swimtime="00:02:21.76" lane="3" heatid="52003" points="344">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:07.44" />
                    <SPLIT distance="150" swimtime="00:01:45.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="786" eventid="42" swimtime="00:00:30.43" lane="2" heatid="42004" points="365" />
                <RESULT resultid="787" eventid="32" swimtime="00:01:01.79" lane="4" heatid="32007" points="382">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172" birthdate="2008-01-01" gender="F" lastname="Johannsohn" firstname="Zoe Tabea" license="390534" nation="GER">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:36.33" heatid="27009" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:13.61" heatid="33009" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:32.87" heatid="41011" lane="3" />
                <ENTRY eventid="45" entrytime="00:01:21.50" heatid="45007" lane="1" />
                <ENTRY eventid="53" entrytime="00:02:43.15" heatid="53003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="788" eventid="27" swimtime="00:00:36.46" lane="3" heatid="27009" points="471" />
                <RESULT resultid="789" eventid="33" swimtime="00:01:14.23" lane="3" heatid="33009" points="441">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="790" eventid="41" swimtime="00:00:33.71" lane="3" heatid="41011" points="378" />
                <RESULT resultid="791" eventid="45" swimtime="00:01:22.78" lane="1" heatid="45007" points="427">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="792" eventid="53" swimtime="00:02:46.04" lane="4" heatid="53003" points="395">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:02:04.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173" birthdate="2003-01-01" gender="M" lastname="Josefus" firstname="Sören" license="294790">
              <ENTRIES>
                <ENTRY eventid="30" entrytime="00:01:01.48" heatid="30003" lane="2" />
                <ENTRY eventid="52" entrytime="00:02:10.67" heatid="52005" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:27.07" heatid="42008" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="793" eventid="30" swimtime="00:01:01.92" lane="2" heatid="30003" points="459">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="794" eventid="52" swimtime="00:02:08.21" lane="4" heatid="52005" points="465">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                    <SPLIT distance="100" swimtime="00:01:03.61" />
                    <SPLIT distance="150" swimtime="00:01:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="795" eventid="42" swimtime="00:00:27.65" lane="3" heatid="42008" points="486" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="174" birthdate="2008-01-01" gender="M" lastname="Kult" firstname="Lenn" license="365315">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.54" heatid="44008" lane="3" />
                <ENTRY eventid="48" entrytime="00:01:13.67" heatid="48002" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:33.21" heatid="26004" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:01.12" heatid="32006" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="796" eventid="44" swimtime="00:00:27.73" lane="3" heatid="44008" points="384" />
                <RESULT resultid="797" eventid="48" swimtime="00:01:13.11" lane="2" heatid="48002" points="288">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="798" eventid="26" swimtime="00:00:33.39" lane="4" heatid="26004" points="290" />
                <RESULT resultid="799" eventid="32" swimtime="00:01:02.05" lane="2" heatid="32006" points="377">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="175" birthdate="2012-01-01" gender="M" lastname="Li" firstname="Joshua" license="437425" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:07.06" heatid="2006" lane="2" />
                <ENTRY eventid="6" entrytime="00:01:16.88" heatid="6012" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:34.11" heatid="18015" lane="2" />
                <ENTRY eventid="22" entrytime="00:02:29.82" heatid="22005" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="800" eventid="2" swimtime="00:01:08.19" lane="2" heatid="2006" points="344">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="801" eventid="6" swimtime="00:01:17.28" lane="2" heatid="6012" points="366">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="802" eventid="18" swimtime="00:00:34.89" lane="2" heatid="18015" points="365" />
                <RESULT resultid="803" eventid="22" swimtime="00:02:30.35" lane="2" heatid="22005" points="387">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:12.91" />
                    <SPLIT distance="150" swimtime="00:01:56.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="176" birthdate="2006-01-01" gender="M" lastname="Littmann" firstname="Finn" license="345608" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.60" heatid="44013" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:03.30" heatid="34005" lane="3" />
                <ENTRY eventid="32" entrytime="00:00:55.06" heatid="32013" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="804" eventid="44" swimtime="00:00:24.26" lane="1" heatid="44013" points="573" />
                <RESULT resultid="805" eventid="34" swimtime="00:01:01.52" lane="3" heatid="34005" points="513">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="806" eventid="32" swimtime="00:00:53.49" lane="4" heatid="32013" points="589">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="177" birthdate="2006-01-01" gender="M" lastname="Mehnert" firstname="Patrick" license="341888">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:29.40" heatid="28011" lane="2" />
                <ENTRY eventid="30" entrytime="00:01:01.25" heatid="30006" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:05.50" heatid="46007" lane="2" />
                <ENTRY eventid="62" entrytime="00:00:29.30" heatid="62001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="807" eventid="28" swimtime="00:00:29.30" lane="2" heatid="28011" points="617" />
                <RESULT resultid="808" eventid="30" status="DNS" swimtime="00:00:00.00" lane="4" heatid="30006" />
                <RESULT resultid="809" eventid="46" swimtime="00:01:05.01" lane="2" heatid="46007" points="614">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2327" eventid="62" swimtime="00:00:29.07" lane="2" heatid="62001" points="632" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="178" birthdate="2010-01-01" gender="M" lastname="Pilz" firstname="Arvid" license="410264" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.38" heatid="44009" lane="3" />
                <ENTRY eventid="30" entrytime="00:01:05.71" heatid="30002" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:29.10" heatid="42006" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:01.60" heatid="32006" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="810" eventid="44" swimtime="00:00:27.30" lane="3" heatid="44009" points="402" />
                <RESULT resultid="811" eventid="30" swimtime="00:01:04.20" lane="2" heatid="30002" points="412">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="812" eventid="42" swimtime="00:00:28.80" lane="4" heatid="42006" points="430" />
                <RESULT resultid="813" eventid="32" swimtime="00:01:01.45" lane="1" heatid="32006" points="388">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="179" birthdate="2010-01-01" gender="M" lastname="Richter" firstname="Toni" license="415137" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:29.02" heatid="44005" lane="2" />
                <ENTRY eventid="52" entrytime="00:02:33.29" heatid="52003" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:31.76" heatid="42004" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:04.79" heatid="32004" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="814" eventid="44" swimtime="00:00:28.58" lane="2" heatid="44005" points="350" />
                <RESULT resultid="815" eventid="52" swimtime="00:02:30.97" lane="4" heatid="52003" points="285">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="816" eventid="42" swimtime="00:00:31.27" lane="1" heatid="42004" points="336" />
                <RESULT resultid="817" eventid="32" swimtime="00:01:04.71" lane="2" heatid="32004" points="332">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="180" birthdate="2008-01-01" gender="F" lastname="Schreiber" firstname="Gretha" license="365675">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:28.68" heatid="43013" lane="2" />
                <ENTRY eventid="51" entrytime="00:02:19.84" heatid="51002" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:02.16" heatid="31012" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="818" eventid="43" swimtime="00:00:28.88" lane="2" heatid="43013" points="500" />
                <RESULT resultid="819" eventid="51" swimtime="00:02:21.02" lane="2" heatid="51002" points="478">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:06.72" />
                    <SPLIT distance="150" swimtime="00:01:44.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="820" eventid="31" swimtime="00:01:04.42" lane="3" heatid="31012" points="474">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="181" birthdate="2011-01-01" gender="F" lastname="Türk" firstname="Emilia" license="408039" nation="GER">
              <ENTRIES>
                <ENTRY eventid="47" entrytime="00:01:17.06" heatid="47005" lane="2" />
                <ENTRY eventid="51" entrytime="00:02:30.49" heatid="51000" lane="0" />
                <ENTRY eventid="25" entrytime="00:00:36.26" heatid="25006" lane="3" />
                <ENTRY eventid="35" entrytime="00:02:44.97" heatid="35003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="821" eventid="47" status="WDR" swimtime="00:00:00.00" lane="2" heatid="47005" />
                <RESULT resultid="822" eventid="51" status="WDR" swimtime="00:00:00.00" lane="0" heatid="51000" />
                <RESULT resultid="823" eventid="25" status="WDR" swimtime="00:00:00.00" lane="3" heatid="25006" />
                <RESULT resultid="824" eventid="35" status="WDR" swimtime="00:00:00.00" lane="4" heatid="35003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182" birthdate="2008-01-01" gender="M" lastname="Uhlig" firstname="Florian" license="368939" nation="GER">
              <ENTRIES>
                <ENTRY eventid="46" entrytime="00:01:24.00" heatid="46002" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:08.16" heatid="32004" lane="3" />
                <ENTRY eventid="36" entrytime="00:02:57.63" heatid="36001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="825" eventid="46" swimtime="00:01:32.06" lane="1" heatid="46002" points="216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="826" eventid="32" swimtime="00:01:07.32" lane="3" heatid="32004" points="295">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="827" eventid="36" swimtime="00:02:58.08" lane="2" heatid="36001" points="208">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:28.07" />
                    <SPLIT distance="150" swimtime="00:02:14.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183" birthdate="2010-01-01" gender="F" lastname="Uhlig" firstname="Julia" license="410268">
              <ENTRIES>
                <ENTRY eventid="25" entrytime="00:00:36.32" heatid="25003" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:11.87" heatid="31006" lane="4" />
                <ENTRY eventid="35" entrytime="00:02:54.31" heatid="35002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="828" eventid="25" status="DNS" swimtime="00:00:00.00" lane="1" heatid="25003" />
                <RESULT resultid="829" eventid="31" status="DNS" swimtime="00:00:00.00" lane="4" heatid="31006" />
                <RESULT resultid="830" eventid="35" status="DNS" swimtime="00:00:00.00" lane="4" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="184" birthdate="2010-01-01" gender="F" lastname="Zeiger" firstname="Hanna" license="410273">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:29.98" heatid="43008" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:36.64" heatid="27008" lane="4" />
                <ENTRY eventid="45" entrytime="00:01:21.38" heatid="45006" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="831" eventid="43" swimtime="00:00:30.00" lane="1" heatid="43008" points="446" />
                <RESULT resultid="832" eventid="27" swimtime="00:00:37.57" lane="4" heatid="27008" points="430" />
                <RESULT resultid="833" eventid="45" swimtime="00:01:21.79" lane="3" heatid="45006" points="443">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:42.25" lane="4" heatid="40003" />
                <ENTRY eventid="72" entrytime="00:01:51.52" lane="4" heatid="72003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="762" eventid="40" swimtime="00:01:39.35" lane="4" heatid="40003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                    <SPLIT distance="100" swimtime="00:00:49.75" />
                    <SPLIT distance="150" swimtime="00:01:15.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="169" number="1" />
                    <RELAYPOSITION athleteid="177" number="2" />
                    <RELAYPOSITION athleteid="173" number="3" />
                    <RELAYPOSITION athleteid="176" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="763" eventid="72" swimtime="00:01:48.90" lane="4" heatid="72003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:00:57.93" />
                    <SPLIT distance="150" swimtime="00:01:25.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="173" number="1" />
                    <RELAYPOSITION athleteid="177" number="2" />
                    <RELAYPOSITION athleteid="169" number="3" />
                    <RELAYPOSITION athleteid="176" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:01:59.67" lane="3" heatid="39002" />
                <ENTRY eventid="71" entrytime="00:02:10.00" lane="3" heatid="71003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="764" eventid="39" swimtime="00:01:58.04" lane="3" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                    <SPLIT distance="100" swimtime="00:00:58.38" />
                    <SPLIT distance="150" swimtime="00:01:28.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="184" number="1" />
                    <RELAYPOSITION athleteid="180" number="2" />
                    <RELAYPOSITION athleteid="167" number="3" />
                    <RELAYPOSITION athleteid="172" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="765" eventid="71" swimtime="00:02:10.57" lane="3" heatid="71003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:01:09.26" />
                    <SPLIT distance="150" swimtime="00:01:41.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="180" number="1" />
                    <RELAYPOSITION athleteid="184" number="2" />
                    <RELAYPOSITION athleteid="172" number="3" />
                    <RELAYPOSITION athleteid="167" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC Eintracht Berlin e.V." nation="GER" region="3" code="5673">
          <ATHLETES>
            <ATHLETE athleteid="133" birthdate="2010-01-01" gender="F" lastname="Brömme" firstname="Lana Marie" license="441656" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:37.22" heatid="43002" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:28.67" heatid="47002" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:30.00" heatid="33002" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:40.28" heatid="41002" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:40.79" heatid="25002" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:23.08" heatid="31002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="611" eventid="43" swimtime="00:00:36.73" lane="3" heatid="43002" points="243" />
                <RESULT resultid="612" eventid="47" status="DSQ" swimtime="00:01:33.95" lane="4" heatid="47002" comment="Bei der ersten Wende wurde die Wand nicht berührt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="613" eventid="33" swimtime="00:01:33.25" lane="3" heatid="33002" points="222">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="614" eventid="41" swimtime="00:00:42.05" lane="3" heatid="41002" points="194" />
                <RESULT resultid="615" eventid="25" swimtime="00:00:41.99" lane="1" heatid="25002" points="217" />
                <RESULT resultid="616" eventid="31" swimtime="00:01:26.63" lane="1" heatid="31002" points="195">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="134" birthdate="2009-01-01" gender="F" lastname="Cappelli" firstname="Emma" license="386111" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:29.45" heatid="43009" lane="4" />
                <ENTRY eventid="29" entrytime="00:01:12.80" heatid="29005" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:32.55" heatid="41006" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:07.15" heatid="31008" lane="1" />
                <ENTRY eventid="63" entrytime="00:00:31.75" heatid="63001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="617" eventid="43" swimtime="00:00:29.57" lane="4" heatid="43009" points="466" />
                <RESULT resultid="618" eventid="29" swimtime="00:01:13.15" lane="1" heatid="29005" points="403">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="619" eventid="41" swimtime="00:00:31.75" lane="3" heatid="41006" points="452" />
                <RESULT resultid="620" eventid="31" swimtime="00:01:06.30" lane="1" heatid="31008" points="435">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2334" eventid="63" swimtime="00:00:31.47" lane="4" heatid="63001" points="464" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="135" birthdate="2010-01-01" gender="F" lastname="Dorn" firstname="Anne" license="435621" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:31.60" heatid="43006" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:41.18" heatid="27004" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:38.02" heatid="41004" lane="3" />
                <ENTRY eventid="45" entrytime="00:01:31.61" heatid="45003" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:13.92" heatid="31005" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="621" eventid="43" swimtime="00:00:30.19" lane="2" heatid="43006" points="438" />
                <RESULT resultid="622" eventid="27" swimtime="00:00:39.18" lane="3" heatid="27004" points="379" />
                <RESULT resultid="623" eventid="41" swimtime="00:00:36.53" lane="3" heatid="41004" points="297" />
                <RESULT resultid="624" eventid="45" swimtime="00:01:30.39" lane="2" heatid="45003" points="328">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="625" eventid="31" swimtime="00:01:10.72" lane="1" heatid="31005" points="358">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="136" birthdate="2011-01-01" gender="M" lastname="Feige" firstname="Bennet" license="441662" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:30.00" heatid="44004" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:41.29" heatid="28002" lane="2" />
                <ENTRY eventid="34" entrytime="00:01:21.70" heatid="34002" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:36.33" heatid="42003" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:37.14" heatid="26003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="626" eventid="44" swimtime="00:00:31.01" lane="3" heatid="44004" points="274" />
                <RESULT resultid="627" eventid="28" status="DSQ" swimtime="00:00:40.24" lane="2" heatid="28002" comment="Beim Zielanschlag hat der Sportler nicht mit beiden Händen gleichzeitig angeschlagen." />
                <RESULT resultid="628" eventid="34" swimtime="00:01:18.57" lane="2" heatid="34002" points="246">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="629" eventid="42" swimtime="00:00:34.00" lane="4" heatid="42003" points="261" />
                <RESULT resultid="630" eventid="26" swimtime="00:00:36.11" lane="4" heatid="26003" points="229" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="137" birthdate="2009-01-01" gender="M" lastname="Kohl" firstname="Roman" license="463367" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:30.00" heatid="44004" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:41.87" heatid="28002" lane="3" />
                <ENTRY eventid="34" entrytime="00:01:23.29" heatid="34002" lane="3" />
                <ENTRY eventid="52" entrytime="00:02:40.00" heatid="52002" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:36.29" heatid="42003" lane="1" />
                <ENTRY eventid="54" entrytime="00:03:03.31" heatid="54001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="631" eventid="44" swimtime="00:00:29.80" lane="2" heatid="44004" points="309" />
                <RESULT resultid="632" eventid="28" swimtime="00:00:39.18" lane="3" heatid="28002" points="258" />
                <RESULT resultid="633" eventid="34" swimtime="00:01:20.52" lane="3" heatid="34002" points="229">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="634" eventid="52" swimtime="00:02:33.96" lane="2" heatid="52002" points="268">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                    <SPLIT distance="150" swimtime="00:01:55.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="635" eventid="42" swimtime="00:00:34.51" lane="1" heatid="42003" points="250" />
                <RESULT resultid="636" eventid="54" status="DSQ" swimtime="00:02:55.86" lane="2" heatid="54001" comment="Vor der zweiten Wende wurde ein Brustarmzug durchgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:26.90" />
                    <SPLIT distance="150" swimtime="00:02:17.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="138" birthdate="2011-01-01" gender="F" lastname="Krüger" firstname="Emilia" license="428927" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:34.66" heatid="43003" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:43.34" heatid="27003" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:27.38" heatid="33003" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:39.21" heatid="41003" lane="3" />
                <ENTRY eventid="45" entrytime="00:01:36.23" heatid="45002" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:18.30" heatid="31003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="637" eventid="43" swimtime="00:00:35.38" lane="2" heatid="43003" points="272" />
                <RESULT resultid="638" eventid="27" swimtime="00:00:43.50" lane="2" heatid="27003" points="277" />
                <RESULT resultid="639" eventid="33" swimtime="00:01:29.07" lane="2" heatid="33003" points="255">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="640" eventid="41" swimtime="00:00:39.32" lane="3" heatid="41003" points="238" />
                <RESULT resultid="641" eventid="45" swimtime="00:01:38.46" lane="1" heatid="45002" points="254">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="642" eventid="31" swimtime="00:01:21.62" lane="1" heatid="31003" points="233">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="139" birthdate="1997-01-01" gender="M" lastname="Rodriguez Weber" firstname="Adrian" license="171364" nation="GER">
              <ENTRIES>
                <ENTRY eventid="32" entrytime="00:00:59.99" heatid="32007" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="643" eventid="32" swimtime="00:01:02.48" lane="2" heatid="32007" points="369">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140" birthdate="2010-01-01" gender="F" lastname="Schatalin" firstname="Elena" license="435619" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:29.73" heatid="43008" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:41.03" heatid="27004" lane="2" />
                <ENTRY eventid="47" entrytime="00:01:14.92" heatid="47003" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:34.01" heatid="41005" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:34.41" heatid="25004" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:06.68" heatid="31008" lane="2" />
                <ENTRY eventid="55" entrytime="00:00:34.20" heatid="55001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="644" eventid="43" swimtime="00:00:29.82" lane="3" heatid="43008" points="454" />
                <RESULT resultid="645" eventid="27" swimtime="00:00:39.57" lane="2" heatid="27004" points="368" />
                <RESULT resultid="646" eventid="47" swimtime="00:01:16.27" lane="2" heatid="47003" points="372">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="647" eventid="41" swimtime="00:00:33.59" lane="3" heatid="41005" points="382" />
                <RESULT resultid="648" eventid="25" swimtime="00:00:34.20" lane="3" heatid="25004" points="402" />
                <RESULT resultid="649" eventid="31" swimtime="00:01:07.19" lane="2" heatid="31008" points="418">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2348" eventid="55" swimtime="00:00:33.65" lane="3" heatid="55001" points="422" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="141" birthdate="2009-01-01" gender="M" lastname="Schober" firstname="Florian" license="439713" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.14" heatid="44010" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:32.40" heatid="28009" lane="4" />
                <ENTRY eventid="38" entrytime="00:02:56.35" heatid="38004" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:29.28" heatid="42005" lane="3" />
                <ENTRY eventid="46" entrytime="00:01:13.09" heatid="46003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="650" eventid="44" swimtime="00:00:27.08" lane="1" heatid="44010" points="412" />
                <RESULT resultid="651" eventid="28" swimtime="00:00:33.81" lane="4" heatid="28009" points="401" />
                <RESULT resultid="652" eventid="38" swimtime="00:02:48.53" lane="3" heatid="38004" points="362">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:20.04" />
                    <SPLIT distance="150" swimtime="00:02:06.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="653" eventid="42" swimtime="00:00:30.01" lane="3" heatid="42005" points="380" />
                <RESULT resultid="654" eventid="46" swimtime="00:01:15.95" lane="2" heatid="46003" points="385">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="142" birthdate="2003-01-01" gender="M" lastname="Schulze" firstname="Eric" license="298385" nation="GER">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:31.54" heatid="28011" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:28.00" heatid="42007" lane="2" />
                <ENTRY eventid="46" entrytime="00:01:13.10" heatid="46007" lane="1" />
                <ENTRY eventid="32" entrytime="00:00:59.99" heatid="32008" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="655" eventid="28" swimtime="00:00:32.33" lane="4" heatid="28011" points="459" />
                <RESULT resultid="656" eventid="42" swimtime="00:00:28.39" lane="2" heatid="42007" points="449" />
                <RESULT resultid="657" eventid="46" swimtime="00:01:20.73" lane="1" heatid="46007" points="321">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="658" eventid="32" status="DNS" swimtime="00:00:00.00" lane="3" heatid="32008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143" birthdate="2011-01-01" gender="M" lastname="Sommer" firstname="Erik" license="441664" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:29.44" heatid="44014" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:39.59" heatid="28004" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:16.00" heatid="34006" lane="1" />
                <ENTRY eventid="52" entrytime="00:02:31.34" heatid="52003" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:34.11" heatid="42010" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:04.44" heatid="32010" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="659" eventid="44" swimtime="00:00:28.94" lane="4" heatid="44014" points="338" />
                <RESULT resultid="660" eventid="28" swimtime="00:00:38.59" lane="1" heatid="28004" points="270" />
                <RESULT resultid="661" eventid="34" swimtime="00:01:16.06" lane="1" heatid="34006" points="271">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="662" eventid="52" swimtime="00:02:32.78" lane="1" heatid="52003" points="275">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                    <SPLIT distance="150" swimtime="00:01:51.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="663" eventid="42" swimtime="00:00:32.42" lane="4" heatid="42010" points="301" />
                <RESULT resultid="664" eventid="32" swimtime="00:01:05.39" lane="3" heatid="32010" points="322">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144" birthdate="2007-01-01" gender="M" lastname="Unger" firstname="Tobias" license="404260" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:26.02" heatid="44012" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:28.88" heatid="42006" lane="2" />
                <ENTRY eventid="32" entrytime="00:00:59.99" heatid="32008" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="665" eventid="44" status="WDR" swimtime="00:00:00.00" lane="4" heatid="44012" />
                <RESULT resultid="666" eventid="42" status="WDR" swimtime="00:00:00.00" lane="2" heatid="42006" />
                <RESULT resultid="667" eventid="32" status="WDR" swimtime="00:00:00.00" lane="4" heatid="32008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145" birthdate="2015-01-01" gender="M" lastname="Yuasa" firstname="Jannes Kenji" license="473246" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:47.17" heatid="4013" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:37.88" heatid="10004" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:53.70" heatid="18005" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:31.91" heatid="20008" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="668" eventid="4" swimtime="00:00:41.36" lane="4" heatid="4013" points="152" />
                <RESULT resultid="669" eventid="10" swimtime="00:01:39.73" lane="4" heatid="10004" points="120">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="670" eventid="18" swimtime="00:00:49.59" lane="3" heatid="18005" points="127" />
                <RESULT resultid="671" eventid="20" swimtime="00:01:32.32" lane="1" heatid="20008" points="114">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="146" birthdate="2013-01-01" gender="F" lastname="Yuasa" firstname="Mavie" license="447450" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:37.27" heatid="3023" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:33.29" heatid="7030" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:20.00" heatid="9018" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:35.91" heatid="13016" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:12.80" heatid="19025" lane="3" />
                <ENTRY eventid="35" entrytime="00:03:00.00" heatid="35001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="672" eventid="3" swimtime="00:00:35.88" lane="1" heatid="3023" points="348" />
                <RESULT resultid="673" eventid="7" swimtime="00:00:33.05" lane="1" heatid="7030" points="333" />
                <RESULT resultid="674" eventid="9" swimtime="00:01:23.16" lane="3" heatid="9018" points="313">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="675" eventid="13" swimtime="00:00:34.74" lane="1" heatid="13016" points="345" />
                <RESULT resultid="676" eventid="19" swimtime="00:01:13.17" lane="3" heatid="19025" points="323">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="677" eventid="35" swimtime="00:02:58.56" lane="2" heatid="35001" points="295">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:26.41" />
                    <SPLIT distance="150" swimtime="00:02:12.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147" birthdate="2009-01-01" gender="F" lastname="Zieb" firstname="Anna Florentine" license="405985" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:28.66" heatid="43009" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:35.83" heatid="27008" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:31.35" heatid="41007" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:33.03" heatid="25004" lane="2" />
                <ENTRY eventid="67" entrytime="00:00:28.62" heatid="67001" lane="1" />
                <ENTRY eventid="60" entrytime="00:00:35.74" heatid="60001" lane="4" />
                <ENTRY eventid="55" entrytime="00:00:33.06" heatid="55001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="678" eventid="43" swimtime="00:00:28.62" lane="3" heatid="43009" points="514" />
                <RESULT resultid="679" eventid="27" swimtime="00:00:35.74" lane="1" heatid="27008" points="500" />
                <RESULT resultid="680" eventid="41" swimtime="00:00:32.28" lane="3" heatid="41007" points="430" />
                <RESULT resultid="681" eventid="25" swimtime="00:00:33.06" lane="2" heatid="25004" points="445" />
                <RESULT resultid="2347" eventid="55" swimtime="00:00:32.48" lane="2" heatid="55001" points="469" />
                <RESULT resultid="2322" eventid="60" swimtime="00:00:35.88" lane="4" heatid="60001" points="494" />
                <RESULT resultid="2301" eventid="67" swimtime="00:00:28.75" lane="1" heatid="67001" points="507" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="148" birthdate="2006-01-01" gender="M" lastname="Zieb" firstname="Tom" license="344952" nation="GER">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:33.51" heatid="28006" lane="2" />
                <ENTRY eventid="32" entrytime="00:00:59.99" heatid="32008" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="682" eventid="28" swimtime="00:00:34.26" lane="2" heatid="28006" points="386" />
                <RESULT resultid="683" eventid="32" swimtime="00:01:02.81" lane="1" heatid="32008" points="363">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:44.00" lane="2" heatid="40002" />
                <ENTRY eventid="72" entrytime="00:01:57.07" lane="2" heatid="72002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="606" eventid="40" swimtime="00:01:44.79" lane="2" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                    <SPLIT distance="100" swimtime="00:00:54.38" />
                    <SPLIT distance="150" swimtime="00:01:20.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="141" number="1" />
                    <RELAYPOSITION athleteid="148" number="2" />
                    <RELAYPOSITION athleteid="142" number="3" />
                    <RELAYPOSITION athleteid="139" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="607" eventid="72" swimtime="00:01:57.10" lane="2" heatid="72002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:02.37" />
                    <SPLIT distance="150" swimtime="00:01:29.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="139" number="1" />
                    <RELAYPOSITION athleteid="141" number="2" />
                    <RELAYPOSITION athleteid="142" number="3" />
                    <RELAYPOSITION athleteid="148" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:01:59.00" lane="2" heatid="39002" />
                <ENTRY eventid="71" entrytime="00:02:16.80" lane="1" heatid="71002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="608" eventid="39" swimtime="00:01:58.28" lane="2" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:00:59.89" />
                    <SPLIT distance="150" swimtime="00:01:30.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="134" number="1" />
                    <RELAYPOSITION athleteid="140" number="2" />
                    <RELAYPOSITION athleteid="135" number="3" />
                    <RELAYPOSITION athleteid="147" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="609" eventid="71" swimtime="00:02:16.85" lane="1" heatid="71002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:15.05" />
                    <SPLIT distance="150" swimtime="00:01:47.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="140" number="1" />
                    <RELAYPOSITION athleteid="135" number="2" />
                    <RELAYPOSITION athleteid="134" number="3" />
                    <RELAYPOSITION athleteid="147" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:56.50" lane="2" heatid="40001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="610" eventid="40" status="DSQ" swimtime="00:02:04.03" lane="2" heatid="40001" comment="Die Füße des dritten StaffelSportlers hatten den Startblock verlassen, bevor der vorherige StaffelSportler die Wand berührt hatte.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="150" swimtime="00:01:35.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="137" number="1" />
                    <RELAYPOSITION athleteid="145" number="2" />
                    <RELAYPOSITION athleteid="136" number="3" />
                    <RELAYPOSITION athleteid="143" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC Freital" nation="GER" region="12" code="3339">
          <ATHLETES>
            <ATHLETE athleteid="275" birthdate="2013-01-01" gender="F" lastname="Amsel" firstname="Helena" license="448347">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:40.42" heatid="3018" lane="3" />
                <ENTRY eventid="5" entrytime="00:01:34.31" heatid="5015" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:29.63" heatid="9012" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:40.74" heatid="13010" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:43.88" heatid="17020" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1183" eventid="3" swimtime="00:00:41.35" lane="3" heatid="3018" points="227" />
                <RESULT resultid="1184" eventid="5" swimtime="00:01:33.77" lane="1" heatid="5015" points="294">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1185" eventid="9" swimtime="00:01:28.45" lane="1" heatid="9012" points="260">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1186" eventid="13" swimtime="00:00:40.68" lane="2" heatid="13010" points="215" />
                <RESULT resultid="1187" eventid="17" swimtime="00:00:42.14" lane="4" heatid="17020" points="305" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="276" birthdate="2011-01-01" gender="M" lastname="Börner" firstname="Fynn" license="425572">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:34.77" heatid="28008" lane="2" />
                <ENTRY eventid="34" entrytime="00:01:12.28" heatid="34006" lane="2" />
                <ENTRY eventid="38" entrytime="00:02:53.78" heatid="38004" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:34.76" heatid="26007" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:08.84" heatid="32004" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1188" eventid="28" swimtime="00:00:34.84" lane="2" heatid="28008" points="367" />
                <RESULT resultid="1189" eventid="34" swimtime="00:01:12.71" lane="2" heatid="34006" points="311">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1190" eventid="38" swimtime="00:02:52.87" lane="2" heatid="38004" points="335">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:23.80" />
                    <SPLIT distance="150" swimtime="00:02:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1191" eventid="26" swimtime="00:00:34.17" lane="1" heatid="26007" points="270" />
                <RESULT resultid="1192" eventid="32" swimtime="00:01:06.60" lane="4" heatid="32004" points="305">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="277" birthdate="2010-01-01" gender="F" lastname="Gahner" firstname="Masine" license="406268">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:29.00" heatid="43009" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:37.77" heatid="27005" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:12.86" heatid="33008" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:31.59" heatid="41007" lane="1" />
                <ENTRY eventid="45" entrytime="00:01:27.08" heatid="45006" lane="4" />
                <ENTRY eventid="67" entrytime="00:00:28.59" heatid="67001" lane="3" />
                <ENTRY eventid="59" entrytime="00:00:37.41" heatid="59001" lane="4" />
                <ENTRY eventid="63" entrytime="00:00:31.52" heatid="63001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1193" eventid="43" swimtime="00:00:28.59" lane="1" heatid="43009" points="515" />
                <RESULT resultid="1194" eventid="27" swimtime="00:00:37.41" lane="3" heatid="27005" points="436" />
                <RESULT resultid="1195" eventid="33" swimtime="00:01:11.90" lane="4" heatid="33008" points="485">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1196" eventid="41" swimtime="00:00:31.52" lane="1" heatid="41007" points="462" />
                <RESULT resultid="1197" eventid="45" swimtime="00:01:23.14" lane="4" heatid="45006" points="421">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2318" eventid="59" swimtime="00:00:37.59" lane="4" heatid="59001" points="429" />
                <RESULT resultid="2333" eventid="63" swimtime="00:00:31.09" lane="1" heatid="63001" points="482" />
                <RESULT resultid="2300" eventid="67" swimtime="00:00:28.81" lane="3" heatid="67001" points="504" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="278" birthdate="2011-01-01" gender="M" lastname="Hentsch" firstname="Oskar René" license="425566">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:42.29" heatid="28002" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:19.96" heatid="34003" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:37.70" heatid="42002" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:36.73" heatid="26003" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:11.89" heatid="32003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1198" eventid="28" swimtime="00:00:42.58" lane="1" heatid="28002" points="201" />
                <RESULT resultid="1199" eventid="34" swimtime="00:01:20.42" lane="1" heatid="34003" points="230">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1200" eventid="42" swimtime="00:00:36.69" lane="3" heatid="42002" points="208" />
                <RESULT resultid="1201" eventid="26" swimtime="00:00:36.78" lane="1" heatid="26003" points="217" />
                <RESULT resultid="1202" eventid="32" swimtime="00:01:10.79" lane="1" heatid="32003" points="254">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="279" birthdate="2010-01-01" gender="F" lastname="Heuer" firstname="Lia-Kiara" license="413355">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.16" heatid="43008" lane="4" />
                <ENTRY eventid="29" entrytime="00:01:19.02" heatid="29005" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:15.37" heatid="33005" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:33.95" heatid="41005" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:07.33" heatid="31008" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1203" eventid="43" swimtime="00:00:30.21" lane="4" heatid="43008" points="437" />
                <RESULT resultid="1204" eventid="29" swimtime="00:01:21.13" lane="4" heatid="29005" points="295">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1205" eventid="33" status="DNS" swimtime="00:00:00.00" lane="4" heatid="33005" />
                <RESULT resultid="1206" eventid="41" swimtime="00:00:34.02" lane="2" heatid="41005" points="368" />
                <RESULT resultid="1207" eventid="31" swimtime="00:01:09.60" lane="4" heatid="31008" points="376">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="280" birthdate="2012-01-01" gender="M" lastname="Kretzschmar" firstname="Nils" license="438792">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:34.91" heatid="2006" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:27.96" heatid="8025" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:34.62" heatid="14012" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:37.84" heatid="18015" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:06.01" heatid="20022" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1208" eventid="2" swimtime="00:01:26.96" lane="4" heatid="2006" points="165">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1209" eventid="8" swimtime="00:00:28.03" lane="2" heatid="8025" points="372" />
                <RESULT resultid="1210" eventid="14" swimtime="00:00:33.82" lane="4" heatid="14012" points="265" />
                <RESULT resultid="1211" eventid="18" swimtime="00:00:37.98" lane="1" heatid="18015" points="283" />
                <RESULT resultid="1212" eventid="20" swimtime="00:01:05.83" lane="3" heatid="20022" points="316">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="281" birthdate="2011-01-01" gender="M" lastname="Kupske" firstname="Julien" license="425568">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:29.09" heatid="44014" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:36.50" heatid="28008" lane="3" />
                <ENTRY eventid="34" entrytime="00:01:14.29" heatid="34006" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:33.98" heatid="42010" lane="1" />
                <ENTRY eventid="46" entrytime="00:01:23.51" heatid="46004" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1213" eventid="44" swimtime="00:00:28.20" lane="2" heatid="44014" points="365" />
                <RESULT resultid="1214" eventid="28" swimtime="00:00:37.84" lane="3" heatid="28008" points="286" />
                <RESULT resultid="1215" eventid="34" swimtime="00:01:14.73" lane="3" heatid="34006" points="286">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1216" eventid="42" swimtime="00:00:32.58" lane="1" heatid="42010" points="297" />
                <RESULT resultid="1217" eventid="46" swimtime="00:01:24.85" lane="3" heatid="46004" points="276">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="282" birthdate="2013-01-01" gender="M" lastname="Lehmann" firstname="Nicklas" license="447310">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:39.88" heatid="2001" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:30.10" heatid="8024" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:34.52" heatid="14011" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:39.62" heatid="18014" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:12.63" heatid="20016" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1218" eventid="2" swimtime="00:01:22.27" lane="2" heatid="2001" points="195">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1219" eventid="8" swimtime="00:00:28.84" lane="3" heatid="8024" points="341" />
                <RESULT resultid="1220" eventid="14" swimtime="00:00:32.63" lane="1" heatid="14011" points="296" />
                <RESULT resultid="1221" eventid="18" swimtime="00:00:39.51" lane="3" heatid="18014" points="251" />
                <RESULT resultid="1222" eventid="20" swimtime="00:01:09.71" lane="3" heatid="20016" points="266">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="283" birthdate="2009-01-01" gender="F" lastname="Lorenz" firstname="Sophia" license="402585">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.43" heatid="43007" lane="2" />
                <ENTRY eventid="47" entrytime="00:01:17.49" heatid="47003" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:33.71" heatid="41006" lane="1" />
                <ENTRY eventid="25" entrytime="00:00:35.56" heatid="25003" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:07.10" heatid="31008" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1223" eventid="43" swimtime="00:00:30.68" lane="2" heatid="43007" points="417" />
                <RESULT resultid="1224" eventid="47" swimtime="00:01:19.80" lane="1" heatid="47003" points="325">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1225" eventid="41" swimtime="00:00:35.37" lane="1" heatid="41006" points="327" />
                <RESULT resultid="1226" eventid="25" swimtime="00:00:36.76" lane="2" heatid="25003" points="324" />
                <RESULT resultid="1227" eventid="31" swimtime="00:01:13.01" lane="3" heatid="31008" points="326">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="284" birthdate="2013-01-01" gender="F" lastname="Mäke" firstname="Elsa" license="448348">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:38.23" heatid="3023" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:34.71" heatid="7024" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:28.10" heatid="9012" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:22.82" heatid="15019" lane="1" />
                <ENTRY eventid="21" entrytime="00:03:09.47" heatid="21003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1228" eventid="3" swimtime="00:00:38.00" lane="4" heatid="3023" points="293" />
                <RESULT resultid="1229" eventid="7" swimtime="00:00:34.05" lane="3" heatid="7024" points="305" />
                <RESULT resultid="1230" eventid="9" swimtime="00:01:25.95" lane="3" heatid="9012" points="284">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1231" eventid="15" swimtime="00:01:23.32" lane="1" heatid="15019" points="285">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1232" eventid="21" swimtime="00:03:05.07" lane="2" heatid="21003" points="285">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                    <SPLIT distance="100" swimtime="00:01:26.03" />
                    <SPLIT distance="150" swimtime="00:02:22.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="285" birthdate="2010-01-01" gender="F" lastname="Mann" firstname="Emma" license="418262">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:34.30" heatid="43004" lane="1" />
                <ENTRY eventid="29" entrytime="00:01:30.73" heatid="29001" lane="1" />
                <ENTRY eventid="33" entrytime="00:01:28.91" heatid="33003" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:38.53" heatid="41004" lane="4" />
                <ENTRY eventid="45" entrytime="00:01:35.01" heatid="45002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1233" eventid="43" swimtime="00:00:33.79" lane="1" heatid="43004" points="312" />
                <RESULT resultid="1234" eventid="29" swimtime="00:01:39.38" lane="1" heatid="29001" points="160">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1235" eventid="33" swimtime="00:01:26.55" lane="3" heatid="33003" points="278">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1236" eventid="41" swimtime="00:00:40.12" lane="4" heatid="41004" points="224" />
                <RESULT resultid="1237" eventid="45" swimtime="00:01:36.83" lane="2" heatid="45002" points="267">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="286" birthdate="2010-01-01" gender="M" lastname="Neubert" firstname="Lino" license="413354">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:31.40" heatid="44003" lane="2" />
                <ENTRY eventid="48" entrytime="00:01:22.90" heatid="48001" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:37.63" heatid="42002" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:37.85" heatid="26002" lane="3" />
                <ENTRY eventid="32" entrytime="00:01:11.79" heatid="32003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1238" eventid="44" swimtime="00:00:31.94" lane="2" heatid="44003" points="251" />
                <RESULT resultid="1239" eventid="48" swimtime="00:01:18.98" lane="2" heatid="48001" points="229">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1240" eventid="42" swimtime="00:00:37.54" lane="2" heatid="42002" points="194" />
                <RESULT resultid="1241" eventid="26" swimtime="00:00:37.09" lane="3" heatid="26002" points="211" />
                <RESULT resultid="1242" eventid="32" swimtime="00:01:12.08" lane="3" heatid="32003" points="240">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="287" birthdate="2011-01-01" gender="F" lastname="Neumann" firstname="Antonia" license="429632">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:31.28" heatid="43011" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:37.62" heatid="27007" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:18.47" heatid="33007" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:35.68" heatid="25006" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:25.53" heatid="45005" lane="2" />
                <ENTRY eventid="59" entrytime="00:00:37.06" heatid="59001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1243" eventid="43" swimtime="00:00:30.25" lane="4" heatid="43011" points="435" />
                <RESULT resultid="1244" eventid="27" swimtime="00:00:37.06" lane="2" heatid="27007" points="448" />
                <RESULT resultid="1245" eventid="33" swimtime="00:01:18.21" lane="3" heatid="33007" points="377">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1246" eventid="25" swimtime="00:00:35.58" lane="2" heatid="25006" points="357" />
                <RESULT resultid="1247" eventid="45" swimtime="00:01:25.05" lane="2" heatid="45005" points="394">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2317" eventid="59" swimtime="00:00:37.05" lane="1" heatid="59001" points="448" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="288" birthdate="2010-01-01" gender="M" lastname="Pink" firstname="Adrian" license="413359">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:28.48" heatid="44006" lane="3" />
                <ENTRY eventid="30" entrytime="00:01:18.52" heatid="30001" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:13.63" heatid="34004" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:32.92" heatid="26004" lane="3" />
                <ENTRY eventid="32" entrytime="00:01:02.73" heatid="32005" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1248" eventid="44" swimtime="00:00:27.75" lane="3" heatid="44006" points="383" />
                <RESULT resultid="1249" eventid="30" swimtime="00:01:15.39" lane="1" heatid="30001" points="254">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1250" eventid="34" swimtime="00:01:12.50" lane="2" heatid="34004" points="314">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1251" eventid="26" swimtime="00:00:32.12" lane="3" heatid="26004" points="326" />
                <RESULT resultid="1252" eventid="32" swimtime="00:01:02.69" lane="3" heatid="32005" points="365">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="289" birthdate="2010-01-01" gender="F" lastname="Röder" firstname="Pauline" license="406267">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:34.60" heatid="43004" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:44.36" heatid="27002" lane="2" />
                <ENTRY eventid="47" entrytime="00:01:26.27" heatid="47002" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:36.75" heatid="41004" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:35.13" heatid="45002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1253" eventid="43" swimtime="00:00:34.45" lane="4" heatid="43004" points="294" />
                <RESULT resultid="1254" eventid="27" swimtime="00:00:43.66" lane="2" heatid="27002" points="274" />
                <RESULT resultid="1255" eventid="47" swimtime="00:01:27.36" lane="1" heatid="47002" points="248">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1256" eventid="41" swimtime="00:00:36.24" lane="2" heatid="41004" points="304" />
                <RESULT resultid="1257" eventid="45" swimtime="00:01:36.45" lane="3" heatid="45002" points="270">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="290" birthdate="2007-01-01" gender="M" lastname="Rödig" firstname="Luca Maurice" license="362599">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.45" heatid="44008" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:33.80" heatid="28010" lane="4" />
                <ENTRY eventid="34" entrytime="00:01:09.99" heatid="34008" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:30.32" heatid="42005" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:16.55" heatid="46006" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1258" eventid="44" swimtime="00:00:27.25" lane="2" heatid="44008" points="404" />
                <RESULT resultid="1259" eventid="28" swimtime="00:00:33.43" lane="4" heatid="28010" points="415" />
                <RESULT resultid="1260" eventid="34" status="DNS" swimtime="00:00:00.00" lane="1" heatid="34008" />
                <RESULT resultid="1261" eventid="42" status="DNS" swimtime="00:00:00.00" lane="4" heatid="42005" />
                <RESULT resultid="1262" eventid="46" status="DNS" swimtime="00:00:00.00" lane="4" heatid="46006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="291" birthdate="2009-01-01" gender="F" lastname="Schmidt" firstname="Carolyn" license="385998">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:28.09" heatid="43012" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:38.52" heatid="27005" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:13.40" heatid="33005" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:32.15" heatid="41007" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:02.98" heatid="31011" lane="1" />
                <ENTRY eventid="68" entrytime="00:00:27.88" heatid="68001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1263" eventid="43" swimtime="00:00:27.88" lane="1" heatid="43012" points="556" />
                <RESULT resultid="1264" eventid="27" swimtime="00:00:38.28" lane="4" heatid="27005" points="407" />
                <RESULT resultid="1265" eventid="33" swimtime="00:01:15.09" lane="2" heatid="33005" points="426">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1266" eventid="41" swimtime="00:00:32.16" lane="4" heatid="41007" points="435" />
                <RESULT resultid="1267" eventid="31" swimtime="00:01:02.76" lane="1" heatid="31011" points="513">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2305" eventid="68" swimtime="00:00:27.89" lane="1" heatid="68001" points="555" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="292" birthdate="2006-01-01" gender="M" lastname="Schmidt" firstname="Moritz-Joy" license="347127">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.48" heatid="44013" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:30.57" heatid="28011" lane="3" />
                <ENTRY eventid="34" entrytime="00:00:58.46" heatid="34009" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:25.30" heatid="42013" lane="1" />
                <ENTRY eventid="26" entrytime="00:00:28.54" heatid="26006" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1268" eventid="44" status="DNS" swimtime="00:00:00.00" lane="3" heatid="44013" />
                <RESULT resultid="1269" eventid="28" status="DNS" swimtime="00:00:00.00" lane="3" heatid="28011" />
                <RESULT resultid="1270" eventid="34" status="DNS" swimtime="00:00:00.00" lane="3" heatid="34009" />
                <RESULT resultid="1271" eventid="42" status="DNS" swimtime="00:00:00.00" lane="1" heatid="42013" />
                <RESULT resultid="1272" eventid="26" status="DNS" swimtime="00:00:00.00" lane="3" heatid="26006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="293" birthdate="2011-01-01" gender="M" lastname="Setzer" firstname="Nils" license="425569">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:30.68" heatid="44004" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:39.41" heatid="28008" lane="4" />
                <ENTRY eventid="48" entrytime="00:01:20.00" heatid="48003" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:38.81" heatid="42002" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:09.33" heatid="32003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1273" eventid="44" swimtime="00:00:31.14" lane="1" heatid="44004" points="271" />
                <RESULT resultid="1274" eventid="28" swimtime="00:00:39.00" lane="4" heatid="28008" points="261" />
                <RESULT resultid="1275" eventid="48" swimtime="00:01:21.02" lane="1" heatid="48003" points="212">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1276" eventid="42" swimtime="00:00:38.24" lane="1" heatid="42002" points="184" />
                <RESULT resultid="1277" eventid="32" swimtime="00:01:10.26" lane="2" heatid="32003" points="259">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="294" birthdate="2012-01-01" gender="M" lastname="Wiedmann" firstname="Runar" license="448346">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:08.04" heatid="2006" lane="3" />
                <ENTRY eventid="6" entrytime="00:01:34.68" heatid="6006" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:29.63" heatid="14012" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:44.18" heatid="18009" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:04.48" heatid="20022" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1278" eventid="2" swimtime="00:01:09.96" lane="3" heatid="2006" points="318">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1279" eventid="6" swimtime="00:01:28.69" lane="3" heatid="6006" points="242">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1280" eventid="14" swimtime="00:00:30.80" lane="2" heatid="14012" points="352" />
                <RESULT resultid="1281" eventid="18" swimtime="00:00:40.12" lane="4" heatid="18009" points="240" />
                <RESULT resultid="1282" eventid="20" swimtime="00:01:03.34" lane="2" heatid="20022" points="354">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:01:58.00" lane="3" heatid="39003" />
                <ENTRY eventid="71" entrytime="00:02:12.00" lane="4" heatid="71003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1178" eventid="39" swimtime="00:01:55.19" lane="3" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="100" swimtime="00:00:59.59" />
                    <SPLIT distance="150" swimtime="00:01:27.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="287" number="1" />
                    <RELAYPOSITION athleteid="277" number="2" />
                    <RELAYPOSITION athleteid="279" number="3" />
                    <RELAYPOSITION athleteid="291" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1179" eventid="71" swimtime="00:02:09.78" lane="4" heatid="71003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:11.03" />
                    <SPLIT distance="150" swimtime="00:01:41.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="279" number="1" />
                    <RELAYPOSITION athleteid="287" number="2" />
                    <RELAYPOSITION athleteid="277" number="3" />
                    <RELAYPOSITION athleteid="291" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:50.00" lane="1" heatid="40002" />
                <ENTRY eventid="72" entrytime="00:02:00.00" lane="1" heatid="72002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1180" eventid="40" swimtime="00:01:49.73" lane="1" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.85" />
                    <SPLIT distance="100" swimtime="00:00:53.60" />
                    <SPLIT distance="150" swimtime="00:01:21.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="292" number="1" />
                    <RELAYPOSITION athleteid="281" number="2" />
                    <RELAYPOSITION athleteid="288" number="3" />
                    <RELAYPOSITION athleteid="276" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1181" eventid="72" swimtime="00:02:09.01" lane="1" heatid="72002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:38.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="288" number="1" />
                    <RELAYPOSITION athleteid="276" number="2" />
                    <RELAYPOSITION athleteid="281" number="3" />
                    <RELAYPOSITION athleteid="293" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:00.00" lane="2" heatid="11003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1182" eventid="11" swimtime="00:01:58.33" lane="2" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:01:02.21" />
                    <SPLIT distance="150" swimtime="00:01:30.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="282" number="1" />
                    <RELAYPOSITION athleteid="284" number="2" />
                    <RELAYPOSITION athleteid="294" number="3" />
                    <RELAYPOSITION athleteid="280" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Sportovni klub ASC" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="370" birthdate="2013-01-01" gender="F" lastname="BAKHOUCHE" firstname="Amel" license="0">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:30.90" heatid="5000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:35.03" heatid="7000" lane="0" />
                <ENTRY eventid="9" entrytime="00:01:26.89" heatid="9000" lane="0" />
                <ENTRY eventid="13" entrytime="00:00:41.01" heatid="13000" lane="0" />
                <ENTRY eventid="17" entrytime="00:00:42.60" heatid="17000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:18.86" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1633" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="1634" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="1635" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
                <RESULT resultid="1636" eventid="13" status="WDR" swimtime="00:00:00.00" lane="0" heatid="13000" />
                <RESULT resultid="1637" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
                <RESULT resultid="1638" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="371" birthdate="2013-01-01" gender="F" lastname="BAKHOUCHE" firstname="Safia" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:43.35" heatid="3000" lane="0" />
                <ENTRY eventid="5" entrytime="00:01:40.29" heatid="5000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:35.07" heatid="7000" lane="0" />
                <ENTRY eventid="15" entrytime="00:01:31.90" heatid="15000" lane="0" />
                <ENTRY eventid="17" entrytime="00:00:45.80" heatid="17000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:15.99" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1639" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="1640" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="1641" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="1642" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="1643" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
                <RESULT resultid="1644" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="372" birthdate="2016-01-01" gender="M" lastname="BOUMA" firstname="Sebastián" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:45.10" heatid="4012" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:40.18" heatid="8021" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:36.46" heatid="10009" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:46.77" heatid="14008" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:34.22" heatid="16007" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:24.19" heatid="20018" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1645" eventid="4" swimtime="00:00:44.42" lane="3" heatid="4012" points="123" />
                <RESULT resultid="1646" eventid="8" swimtime="00:00:38.39" lane="4" heatid="8021" points="144" />
                <RESULT resultid="1647" eventid="10" swimtime="00:01:38.50" lane="3" heatid="10009" points="125">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1648" eventid="14" swimtime="00:00:47.45" lane="3" heatid="14008" points="96" />
                <RESULT resultid="1649" eventid="16" swimtime="00:01:37.03" lane="2" heatid="16007" points="123">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1650" eventid="20" swimtime="00:01:29.69" lane="2" heatid="20018" points="124">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="373" birthdate="2015-01-01" gender="F" lastname="CADILOVÁ" firstname="Denisa" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:41.61" heatid="3021" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:34.94" heatid="7028" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:30.14" heatid="9016" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:47.08" heatid="17014" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:17.65" heatid="19023" lane="1" />
                <ENTRY eventid="21" entrytime="00:03:14.31" heatid="21003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1651" eventid="3" swimtime="00:00:40.68" lane="1" heatid="3021" points="239" />
                <RESULT resultid="1652" eventid="7" swimtime="00:00:34.77" lane="3" heatid="7028" points="286" />
                <RESULT resultid="1653" eventid="9" swimtime="00:01:29.33" lane="4" heatid="9016" points="253">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1654" eventid="17" swimtime="00:00:46.07" lane="4" heatid="17014" points="233" />
                <RESULT resultid="1655" eventid="19" swimtime="00:01:16.04" lane="1" heatid="19023" points="288">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1656" eventid="21" swimtime="00:03:14.90" lane="4" heatid="21003" points="244">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                    <SPLIT distance="100" swimtime="00:01:34.07" />
                    <SPLIT distance="150" swimtime="00:02:31.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="374" birthdate="2015-01-01" gender="F" lastname="CAPKOVÁ" firstname="Aneta" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:46.13" heatid="3013" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:40.26" heatid="7016" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:44.84" heatid="9005" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:53.23" heatid="13003" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:43.95" heatid="15008" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:35.39" heatid="19011" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1657" eventid="3" swimtime="00:00:46.09" lane="3" heatid="3013" points="164" />
                <RESULT resultid="1658" eventid="7" swimtime="00:00:39.45" lane="1" heatid="7016" points="196" />
                <RESULT resultid="1659" eventid="9" swimtime="00:01:45.52" lane="3" heatid="9005" points="153">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1660" eventid="13" swimtime="00:00:49.32" lane="4" heatid="13003" points="120" />
                <RESULT resultid="1661" eventid="15" swimtime="00:01:47.43" lane="1" heatid="15008" points="133">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1662" eventid="19" swimtime="00:01:29.86" lane="4" heatid="19011" points="174">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="375" birthdate="2012-01-01" gender="F" lastname="CAPKOVÁ" firstname="Klára" license="0">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:31.88" heatid="43006" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:44.76" heatid="27006" lane="4" />
                <ENTRY eventid="51" entrytime="00:02:41.17" heatid="51001" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:42.44" heatid="41001" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:38.00" heatid="45004" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:13.32" heatid="31005" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1663" eventid="43" swimtime="00:00:33.79" lane="1" heatid="43006" points="312" />
                <RESULT resultid="1664" eventid="27" swimtime="00:00:43.69" lane="4" heatid="27006" points="273" />
                <RESULT resultid="1665" eventid="51" swimtime="00:02:36.76" lane="2" heatid="51001" points="348">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.35" />
                    <SPLIT distance="150" swimtime="00:01:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1666" eventid="41" swimtime="00:00:38.05" lane="2" heatid="41001" points="263" />
                <RESULT resultid="1667" eventid="45" swimtime="00:01:38.32" lane="4" heatid="45004" points="255">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1668" eventid="31" swimtime="00:01:11.79" lane="3" heatid="31005" points="342">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="376" birthdate="2011-01-01" gender="M" lastname="DUFEK" firstname="Matej" license="0">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:29.64" heatid="44005" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:16.62" heatid="34006" lane="4" />
                <ENTRY eventid="52" entrytime="00:02:29.04" heatid="52003" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:33.38" heatid="42010" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:35.73" heatid="26007" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:07.37" heatid="32010" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1669" eventid="44" swimtime="00:00:29.90" lane="1" heatid="44005" points="306" />
                <RESULT resultid="1670" eventid="34" swimtime="00:01:16.08" lane="4" heatid="34006" points="271">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1671" eventid="52" swimtime="00:02:27.21" lane="2" heatid="52003" points="307">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:48.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1672" eventid="42" swimtime="00:00:31.86" lane="3" heatid="42010" points="318" />
                <RESULT resultid="1673" eventid="26" swimtime="00:00:35.35" lane="4" heatid="26007" points="244" />
                <RESULT resultid="1674" eventid="32" swimtime="00:01:04.62" lane="4" heatid="32010" points="334">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="377" birthdate="2015-01-01" gender="F" lastname="ERHARDOVÁ" firstname="Zuzana" license="0">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:43.62" heatid="5009" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:36.88" heatid="7020" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:36.81" heatid="9008" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:46.86" heatid="17014" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:25.36" heatid="19015" lane="1" />
                <ENTRY eventid="21" entrytime="00:03:34.80" heatid="21001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1675" eventid="5" swimtime="00:01:41.94" lane="4" heatid="5009" points="228">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1676" eventid="7" swimtime="00:00:34.16" lane="1" heatid="7020" points="302" />
                <RESULT resultid="1677" eventid="9" swimtime="00:01:33.74" lane="4" heatid="9008" points="219">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1678" eventid="17" swimtime="00:00:47.30" lane="1" heatid="17014" points="215" />
                <RESULT resultid="1679" eventid="19" swimtime="00:01:21.78" lane="1" heatid="19015" points="231">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1680" eventid="21" swimtime="00:03:22.81" lane="1" heatid="21001" points="216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.68" />
                    <SPLIT distance="100" swimtime="00:01:37.09" />
                    <SPLIT distance="150" swimtime="00:02:39.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="378" birthdate="2014-01-01" gender="M" lastname="HAVELKA" firstname="Adam" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:49.71" heatid="4006" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:39.51" heatid="8011" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:40.32" heatid="10003" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:48.47" heatid="14003" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:48.28" heatid="16003" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:28.16" heatid="20009" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1681" eventid="4" status="WDR" swimtime="00:00:00.00" lane="4" heatid="4006" />
                <RESULT resultid="1682" eventid="8" status="WDR" swimtime="00:00:00.00" lane="1" heatid="8011" />
                <RESULT resultid="1683" eventid="10" status="WDR" swimtime="00:00:00.00" lane="1" heatid="10003" />
                <RESULT resultid="1684" eventid="14" status="WDR" swimtime="00:00:00.00" lane="3" heatid="14003" />
                <RESULT resultid="1685" eventid="16" status="WDR" swimtime="00:00:00.00" lane="1" heatid="16003" />
                <RESULT resultid="1686" eventid="20" status="WDR" swimtime="00:00:00.00" lane="4" heatid="20009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="379" birthdate="2009-01-01" gender="M" lastname="JELSA" firstname="Matej" license="0">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:25.83" heatid="44015" lane="1" />
                <ENTRY eventid="30" entrytime="00:01:00.61" heatid="30004" lane="2" />
                <ENTRY eventid="52" entrytime="00:02:07.21" heatid="52005" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:26.83" heatid="42011" lane="2" />
                <ENTRY eventid="32" entrytime="00:00:57.01" heatid="32011" lane="1" />
                <ENTRY eventid="50" entrytime="00:02:17.60" heatid="50002" lane="2" />
                <ENTRY eventid="65" entrytime="00:00:26.89" heatid="65001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1687" eventid="44" swimtime="00:00:26.27" lane="1" heatid="44015" points="451" />
                <RESULT resultid="1688" eventid="30" swimtime="00:01:01.53" lane="2" heatid="30004" points="468">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1689" eventid="52" swimtime="00:02:08.98" lane="3" heatid="52005" points="457">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="100" swimtime="00:01:01.96" />
                    <SPLIT distance="150" swimtime="00:01:35.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1690" eventid="42" swimtime="00:00:26.89" lane="2" heatid="42011" points="529" />
                <RESULT resultid="1691" eventid="32" swimtime="00:00:59.62" lane="1" heatid="32011" points="425">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1692" eventid="50" swimtime="00:02:30.07" lane="2" heatid="50002" points="360">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:51.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2341" eventid="65" swimtime="00:00:26.54" lane="1" heatid="65001" points="550" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="380" birthdate="2014-01-01" gender="M" lastname="JÍLEK" firstname="Tadeás" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:41.74" heatid="4010" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:33.02" heatid="8018" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:25.40" heatid="10000" lane="0" />
                <ENTRY eventid="16" entrytime="00:01:28.59" heatid="16005" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:14.71" heatid="20014" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1693" eventid="4" swimtime="00:00:40.19" lane="1" heatid="4010" points="166" />
                <RESULT resultid="1694" eventid="8" swimtime="00:00:33.98" lane="2" heatid="8018" points="208" />
                <RESULT resultid="1695" eventid="10" status="WDR" swimtime="00:00:00.00" lane="0" heatid="10000" />
                <RESULT resultid="1696" eventid="16" swimtime="00:01:31.65" lane="1" heatid="16005" points="146">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1697" eventid="20" swimtime="00:01:13.85" lane="3" heatid="20014" points="223">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="381" birthdate="2016-01-01" gender="M" lastname="KLIMES" firstname="Viktor" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:02:01.82" heatid="6008" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:41.94" heatid="8008" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:54.83" heatid="18011" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:37.39" heatid="20006" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1698" eventid="6" status="DSQ" swimtime="00:01:54.93" lane="4" heatid="6008" comment="Nach der ersten und dritten Wende hat der Sportler zwei Delphinbeinschläge ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1699" eventid="8" swimtime="00:00:42.37" lane="2" heatid="8008" points="107" />
                <RESULT resultid="1700" eventid="18" swimtime="00:00:55.21" lane="1" heatid="18011" points="92" />
                <RESULT resultid="1701" eventid="20" swimtime="00:01:35.37" lane="4" heatid="20006" points="103">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="382" birthdate="2016-01-01" gender="F" lastname="KNIEZKOVÁ" firstname="Daniela" license="0">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:50.31" heatid="5012" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:43.07" heatid="7012" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:52.53" heatid="17009" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:42.38" heatid="19008" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1702" eventid="5" swimtime="00:01:48.73" lane="1" heatid="5012" points="188">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1703" eventid="7" swimtime="00:00:42.25" lane="1" heatid="7012" points="159" />
                <RESULT resultid="1704" eventid="17" swimtime="00:00:53.04" lane="4" heatid="17009" points="153" />
                <RESULT resultid="1705" eventid="19" swimtime="00:01:37.77" lane="2" heatid="19008" points="135">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="383" birthdate="2007-01-01" gender="F" lastname="KRATOCHVÍLOVÁ" firstname="Monika" license="0">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:33.50" heatid="27009" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:06.59" heatid="33009" lane="2" />
                <ENTRY eventid="37" entrytime="00:02:33.73" heatid="37002" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:11.03" heatid="45007" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:00.24" heatid="31012" lane="2" />
                <ENTRY eventid="53" entrytime="00:02:23.68" heatid="53003" lane="2" />
                <ENTRY eventid="60" entrytime="00:00:34.38" heatid="60001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1706" eventid="27" swimtime="00:00:34.38" lane="2" heatid="27009" points="561" />
                <RESULT resultid="1707" eventid="33" swimtime="00:01:10.38" lane="2" heatid="33009" points="517">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1708" eventid="37" swimtime="00:02:42.01" lane="2" heatid="37002" points="573">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:00.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1709" eventid="45" swimtime="00:01:16.69" lane="2" heatid="45007" points="537">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1710" eventid="31" swimtime="00:01:02.02" lane="2" heatid="31012" points="531">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1711" eventid="53" swimtime="00:02:29.47" lane="2" heatid="53003" points="541">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2321" eventid="60" swimtime="00:00:34.01" lane="1" heatid="60001" points="580" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="384" birthdate="2017-01-01" gender="F" lastname="ORAVCOVÁ" firstname="Alice" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:53.34" heatid="3007" lane="3" />
                <ENTRY eventid="5" entrytime="00:02:23.38" heatid="5002" lane="1" />
                <ENTRY eventid="17" entrytime="00:01:04.35" heatid="17004" lane="4" />
                <ENTRY eventid="19" entrytime="00:02:01.39" heatid="19003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1712" eventid="3" swimtime="00:00:49.65" lane="3" heatid="3007" points="131" />
                <RESULT resultid="1713" eventid="5" swimtime="00:02:11.70" lane="1" heatid="5002" points="106">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1714" eventid="17" swimtime="00:01:03.81" lane="4" heatid="17004" points="87" />
                <RESULT resultid="1715" eventid="19" swimtime="00:01:55.38" lane="1" heatid="19003" points="82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="385" birthdate="2014-01-01" gender="M" lastname="ORAVEC" firstname="Adam" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:52.57" heatid="4003" lane="3" />
                <ENTRY eventid="6" entrytime="00:02:05.89" heatid="6001" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:41.15" heatid="8009" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:43.14" heatid="16003" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:59.95" heatid="18003" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:36.36" heatid="20007" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1716" eventid="4" swimtime="00:00:45.92" lane="3" heatid="4003" points="111" />
                <RESULT resultid="1717" eventid="6" status="DSQ" swimtime="00:02:01.47" lane="3" heatid="6001" comment="Beim Anschlag an der zweiten Wende hat der Sportler nicht mit beiden Händen gleichzeitig angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1718" eventid="8" swimtime="00:00:43.25" lane="2" heatid="8009" points="101" />
                <RESULT resultid="1719" eventid="16" swimtime="00:01:45.33" lane="3" heatid="16003" points="96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1720" eventid="18" swimtime="00:00:56.80" lane="4" heatid="18003" points="84" />
                <RESULT resultid="1721" eventid="20" swimtime="00:01:39.65" lane="4" heatid="20007" points="91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="386" birthdate="2009-01-01" gender="M" lastname="OUREDNÍK" firstname="Adam" license="0">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:25.97" heatid="44015" lane="4" />
                <ENTRY eventid="30" entrytime="00:01:03.02" heatid="30004" lane="1" />
                <ENTRY eventid="52" entrytime="00:02:02.91" heatid="52006" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:28.38" heatid="42011" lane="4" />
                <ENTRY eventid="32" entrytime="00:00:56.52" heatid="32011" lane="3" />
                <ENTRY eventid="50" entrytime="00:02:22.64" heatid="50002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1722" eventid="44" swimtime="00:00:25.87" lane="4" heatid="44015" points="473" />
                <RESULT resultid="1723" eventid="30" swimtime="00:01:03.08" lane="1" heatid="30004" points="434">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1724" eventid="52" swimtime="00:02:04.97" lane="4" heatid="52006" points="502">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="100" swimtime="00:01:01.14" />
                    <SPLIT distance="150" swimtime="00:01:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1725" eventid="42" swimtime="00:00:27.95" lane="4" heatid="42011" points="471" />
                <RESULT resultid="1726" eventid="32" swimtime="00:00:56.01" lane="3" heatid="32011" points="513">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1727" eventid="50" swimtime="00:02:30.73" lane="1" heatid="50002" points="356">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:53.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="387" birthdate="2012-01-01" gender="M" lastname="PAVLÍK" firstname="Marek" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:30.45" heatid="6006" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:33.18" heatid="8018" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:22.37" heatid="10007" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:41.83" heatid="18009" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:15.96" heatid="20014" lane="4" />
                <ENTRY eventid="22" entrytime="00:03:03.33" heatid="22003" lane="2" />
                <ENTRY eventid="38" entrytime="00:03:11.38" heatid="38003" lane="2" />
                <ENTRY eventid="50" entrytime="00:03:43.20" heatid="50000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1728" eventid="6" swimtime="00:01:31.95" lane="2" heatid="6006" points="217">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1729" eventid="8" swimtime="00:00:33.75" lane="1" heatid="8018" points="213" />
                <RESULT resultid="1730" eventid="10" status="DSQ" swimtime="00:01:25.14" lane="2" heatid="10007" comment="Bei der zweiten Wende wurde die Wand nicht berührt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1731" eventid="18" swimtime="00:00:40.48" lane="3" heatid="18009" points="234" />
                <RESULT resultid="1732" eventid="20" swimtime="00:01:14.92" lane="4" heatid="20014" points="214">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1733" eventid="22" swimtime="00:03:01.44" lane="2" heatid="22003" points="220">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:31.02" />
                    <SPLIT distance="150" swimtime="00:02:21.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1734" eventid="38" swimtime="00:03:17.68" lane="2" heatid="38003" points="224">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                    <SPLIT distance="100" swimtime="00:01:35.92" />
                    <SPLIT distance="150" swimtime="00:02:26.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1735" eventid="50" status="WDR" swimtime="00:00:00.00" lane="0" heatid="50000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="388" birthdate="2012-01-01" gender="F" lastname="PAVLÍKOVÁ" firstname="Lucie" license="0">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:31.44" heatid="43010" lane="4" />
                <ENTRY eventid="29" entrytime="00:01:18.54" heatid="29003" lane="4" />
                <ENTRY eventid="47" entrytime="00:01:16.68" heatid="47004" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:35.40" heatid="41008" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:10.30" heatid="31009" lane="4" />
                <ENTRY eventid="35" entrytime="00:02:46.01" heatid="35002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1736" eventid="43" swimtime="00:00:30.89" lane="4" heatid="43010" points="409" />
                <RESULT resultid="1737" eventid="29" swimtime="00:01:18.77" lane="4" heatid="29003" points="323">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1738" eventid="47" swimtime="00:01:15.51" lane="3" heatid="47004" points="384">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1739" eventid="41" swimtime="00:00:33.02" lane="1" heatid="41008" points="402" />
                <RESULT resultid="1740" eventid="31" swimtime="00:01:08.74" lane="4" heatid="31009" points="390">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1741" eventid="35" swimtime="00:02:51.89" lane="1" heatid="35002" points="331">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:02:07.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="389" birthdate="2009-01-01" gender="M" lastname="PAZDÍREK" firstname="Adam" license="0">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.12" heatid="44010" lane="3" />
                <ENTRY eventid="30" entrytime="00:01:04.83" heatid="30003" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:05.91" heatid="34007" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:28.86" heatid="42007" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:14.70" heatid="46003" lane="3" />
                <ENTRY eventid="32" entrytime="00:00:59.00" heatid="32009" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1742" eventid="44" swimtime="00:00:27.49" lane="3" heatid="44010" points="394" />
                <RESULT resultid="1743" eventid="30" swimtime="00:01:07.08" lane="1" heatid="30003" points="361">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1744" eventid="34" swimtime="00:01:13.15" lane="3" heatid="34007" points="305">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1745" eventid="42" swimtime="00:00:30.40" lane="4" heatid="42007" points="366" />
                <RESULT resultid="1746" eventid="46" status="DNS" swimtime="00:00:00.00" lane="3" heatid="46003" />
                <RESULT resultid="1747" eventid="32" swimtime="00:01:01.65" lane="4" heatid="32009" points="384">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="390" birthdate="2015-01-01" gender="M" lastname="PESÁK" firstname="Jan" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:53.83" heatid="6003" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:44.33" heatid="8006" lane="1" />
                <ENTRY eventid="16" entrytime="00:01:57.30" heatid="16002" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:54.62" heatid="18004" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:36.91" heatid="20006" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1748" eventid="6" status="DNS" swimtime="00:00:00.00" lane="3" heatid="6003" />
                <RESULT resultid="1749" eventid="8" status="DNS" swimtime="00:00:00.00" lane="1" heatid="8006" />
                <RESULT resultid="1750" eventid="16" status="DNS" swimtime="00:00:00.00" lane="1" heatid="16002" />
                <RESULT resultid="1751" eventid="18" status="DNS" swimtime="00:00:00.00" lane="2" heatid="18004" />
                <RESULT resultid="1752" eventid="20" status="DNS" swimtime="00:00:00.00" lane="1" heatid="20006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="391" birthdate="2016-01-01" gender="M" lastname="POS" firstname="Antonín" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:02:03.17" heatid="6002" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:58.54" heatid="10001" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:56.00" heatid="18011" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:45.13" heatid="20004" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1753" eventid="6" swimtime="00:02:02.92" lane="3" heatid="6002" points="90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1754" eventid="10" swimtime="00:01:54.95" lane="2" heatid="10001" points="78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1755" eventid="18" swimtime="00:00:56.99" lane="4" heatid="18011" points="83" />
                <RESULT resultid="1756" eventid="20" swimtime="00:01:42.22" lane="4" heatid="20004" points="84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="392" birthdate="2009-01-01" gender="M" lastname="RAK" firstname="Johan" license="0">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.64" heatid="44000" lane="0" />
                <ENTRY eventid="30" entrytime="00:01:16.71" heatid="30000" lane="0" />
                <ENTRY eventid="34" entrytime="00:01:16.94" heatid="34000" lane="0" />
                <ENTRY eventid="42" entrytime="00:00:30.97" heatid="42000" lane="0" />
                <ENTRY eventid="26" entrytime="00:00:35.46" heatid="26000" lane="0" />
                <ENTRY eventid="32" entrytime="00:01:03.31" heatid="32000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1757" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="1758" eventid="30" status="WDR" swimtime="00:00:00.00" lane="0" heatid="30000" />
                <RESULT resultid="1759" eventid="34" status="WDR" swimtime="00:00:00.00" lane="0" heatid="34000" />
                <RESULT resultid="1760" eventid="42" status="WDR" swimtime="00:00:00.00" lane="0" heatid="42000" />
                <RESULT resultid="1761" eventid="26" status="WDR" swimtime="00:00:00.00" lane="0" heatid="26000" />
                <RESULT resultid="1762" eventid="32" status="WDR" swimtime="00:00:00.00" lane="0" heatid="32000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="393" birthdate="2011-01-01" gender="F" lastname="ROUSAROVÁ" firstname="Valentýna" license="0">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:33.91" heatid="43000" lane="0" />
                <ENTRY eventid="47" entrytime="00:01:27.65" heatid="47000" lane="0" />
                <ENTRY eventid="33" entrytime="00:01:28.90" heatid="33000" lane="0" />
                <ENTRY eventid="25" entrytime="00:00:42.16" heatid="25000" lane="0" />
                <ENTRY eventid="31" entrytime="00:01:15.74" heatid="31000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1763" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
                <RESULT resultid="1764" eventid="47" status="WDR" swimtime="00:00:00.00" lane="0" heatid="47000" />
                <RESULT resultid="1765" eventid="33" status="WDR" swimtime="00:00:00.00" lane="0" heatid="33000" />
                <RESULT resultid="1766" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
                <RESULT resultid="1767" eventid="31" status="WDR" swimtime="00:00:00.00" lane="0" heatid="31000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="394" birthdate="2016-01-01" gender="M" lastname="ROZEK" firstname="Michael" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:51.08" heatid="4005" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:48.67" heatid="8004" lane="1" />
                <ENTRY eventid="16" entrytime="00:01:57.08" heatid="16002" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:46.07" heatid="20003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1768" eventid="4" status="DSQ" swimtime="00:00:51.65" lane="4" heatid="4005" comment="Der Sportler hat während der Schwimmstrecke die Rückenlage verlassen." />
                <RESULT resultid="1769" eventid="8" swimtime="00:00:45.51" lane="1" heatid="8004" points="86" />
                <RESULT resultid="1770" eventid="16" swimtime="00:01:56.56" lane="3" heatid="16002" points="71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1771" eventid="20" swimtime="00:01:46.89" lane="2" heatid="20003" points="73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="395" birthdate="2014-01-01" gender="F" lastname="SEBÁNOVÁ" firstname="Linda" license="0">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:30.00" heatid="1002" lane="2" />
                <ENTRY eventid="3" entrytime="00:00:37.80" heatid="3022" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:32.78" heatid="7029" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:37.74" heatid="13011" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:22.94" heatid="15014" lane="3" />
                <ENTRY eventid="21" entrytime="00:03:17.49" heatid="21002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1772" eventid="1" swimtime="00:01:29.31" lane="2" heatid="1002" points="221">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1773" eventid="3" swimtime="00:00:37.76" lane="2" heatid="3022" points="299" />
                <RESULT resultid="1774" eventid="7" swimtime="00:00:32.44" lane="1" heatid="7029" points="353" />
                <RESULT resultid="1775" eventid="13" swimtime="00:00:38.03" lane="2" heatid="13011" points="263" />
                <RESULT resultid="1776" eventid="15" swimtime="00:01:22.00" lane="3" heatid="15014" points="299">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1777" eventid="21" swimtime="00:03:07.70" lane="2" heatid="21002" points="273">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:01:28.15" />
                    <SPLIT distance="150" swimtime="00:02:27.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="396" birthdate="2016-01-01" gender="F" lastname="SIMKOVÁ" firstname="Apollonia" license="0">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:00:50.02" heatid="7007" lane="1" />
                <ENTRY eventid="9" entrytime="00:02:00.52" heatid="9002" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:56.82" heatid="17006" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:48.05" heatid="19005" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1778" eventid="7" swimtime="00:00:47.67" lane="1" heatid="7007" points="111" />
                <RESULT resultid="1779" eventid="9" swimtime="00:02:05.80" lane="3" heatid="9002" points="90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1780" eventid="17" swimtime="00:00:59.07" lane="1" heatid="17006" points="110" />
                <RESULT resultid="1781" eventid="19" swimtime="00:01:52.39" lane="2" heatid="19005" points="89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="397" birthdate="2016-01-01" gender="M" lastname="SINDLÁR" firstname="Benedikt Oliver" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:57.74" heatid="4000" lane="0" />
                <ENTRY eventid="8" entrytime="00:00:44.41" heatid="8000" lane="0" />
                <ENTRY eventid="16" entrytime="00:01:59.79" heatid="16000" lane="0" />
                <ENTRY eventid="20" entrytime="00:01:42.18" heatid="20000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1782" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="1783" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="1784" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="1785" eventid="20" status="WDR" swimtime="00:00:00.00" lane="0" heatid="20000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="398" birthdate="2011-01-01" gender="F" lastname="SKODOVÁ" firstname="Daniela" license="0">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:38.97" heatid="27000" lane="0" />
                <ENTRY eventid="29" entrytime="00:01:15.87" heatid="29000" lane="0" />
                <ENTRY eventid="33" entrytime="00:01:14.74" heatid="33000" lane="0" />
                <ENTRY eventid="41" entrytime="00:00:33.62" heatid="41000" lane="0" />
                <ENTRY eventid="45" entrytime="00:01:22.48" heatid="45000" lane="0" />
                <ENTRY eventid="53" entrytime="00:02:37.70" heatid="53000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1786" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="1787" eventid="29" status="WDR" swimtime="00:00:00.00" lane="0" heatid="29000" />
                <RESULT resultid="1788" eventid="33" status="WDR" swimtime="00:00:00.00" lane="0" heatid="33000" />
                <RESULT resultid="1789" eventid="41" status="WDR" swimtime="00:00:00.00" lane="0" heatid="41000" />
                <RESULT resultid="1790" eventid="45" status="WDR" swimtime="00:00:00.00" lane="0" heatid="45000" />
                <RESULT resultid="1791" eventid="53" status="WDR" swimtime="00:00:00.00" lane="0" heatid="53000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="399" birthdate="2015-01-01" gender="M" lastname="STEHLÍK" firstname="Samuel Patrik" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:33.13" heatid="6009" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:34.70" heatid="8022" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:26.70" heatid="10010" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:42.27" heatid="18012" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:18.12" heatid="20019" lane="3" />
                <ENTRY eventid="22" entrytime="00:03:10.26" heatid="22003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1792" eventid="6" swimtime="00:01:32.12" lane="2" heatid="6009" points="216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1793" eventid="8" swimtime="00:00:35.54" lane="4" heatid="8022" points="182" />
                <RESULT resultid="1794" eventid="10" swimtime="00:01:25.95" lane="3" heatid="10010" points="188">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1795" eventid="18" swimtime="00:00:42.16" lane="2" heatid="18012" points="207" />
                <RESULT resultid="1796" eventid="20" swimtime="00:01:16.30" lane="3" heatid="20019" points="202">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1797" eventid="22" swimtime="00:03:05.66" lane="3" heatid="22003" points="205">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                    <SPLIT distance="100" swimtime="00:01:34.52" />
                    <SPLIT distance="150" swimtime="00:02:24.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="400" birthdate="2012-01-01" gender="F" lastname="STEHLÍKOVÁ" firstname="Linda Wendy" license="0">
              <ENTRIES>
                <ENTRY eventid="29" entrytime="00:01:18.24" heatid="29003" lane="1" />
                <ENTRY eventid="47" entrytime="00:01:15.85" heatid="47004" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:18.19" heatid="33006" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:34.95" heatid="25005" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:10.01" heatid="31009" lane="1" />
                <ENTRY eventid="35" entrytime="00:02:45.34" heatid="35002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1798" eventid="29" swimtime="00:01:18.29" lane="1" heatid="29003" points="329">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1799" eventid="47" swimtime="00:01:15.23" lane="2" heatid="47004" points="388">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1800" eventid="33" swimtime="00:01:18.34" lane="3" heatid="33006" points="375">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1801" eventid="25" swimtime="00:00:35.50" lane="2" heatid="25005" points="359" />
                <RESULT resultid="1802" eventid="31" swimtime="00:01:10.91" lane="1" heatid="31009" points="355">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1803" eventid="35" swimtime="00:02:46.22" lane="2" heatid="35002" points="366">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="150" swimtime="00:02:04.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="401" birthdate="2014-01-01" gender="F" lastname="TANEV" firstname="Emily" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:48.16" heatid="3000" lane="0" />
                <ENTRY eventid="5" entrytime="00:01:55.18" heatid="5000" lane="0" />
                <ENTRY eventid="9" entrytime="00:01:54.41" heatid="9000" lane="0" />
                <ENTRY eventid="15" entrytime="00:01:47.37" heatid="15000" lane="0" />
                <ENTRY eventid="17" entrytime="00:00:54.47" heatid="17000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:41.75" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1804" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="1805" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="1806" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
                <RESULT resultid="1807" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="1808" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
                <RESULT resultid="1809" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="402" birthdate="2016-01-01" gender="F" lastname="TANEV" firstname="Rozálie" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:54.41" heatid="3000" lane="0" />
                <ENTRY eventid="5" entrytime="00:02:11.38" heatid="5000" lane="0" />
                <ENTRY eventid="15" entrytime="00:02:02.86" heatid="15000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:54.93" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1810" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="1811" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="1812" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="1813" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="403" birthdate="2012-01-01" gender="M" lastname="VACA" firstname="Vojtech" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:24.86" heatid="6012" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:30.52" heatid="8025" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:19.47" heatid="10013" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:40.78" heatid="18009" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:06.22" heatid="20022" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1814" eventid="6" swimtime="00:01:24.86" lane="3" heatid="6012" points="276">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1815" eventid="8" swimtime="00:00:29.69" lane="4" heatid="8025" points="313" />
                <RESULT resultid="1816" eventid="10" swimtime="00:01:17.67" lane="4" heatid="10013" points="255">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1817" eventid="18" swimtime="00:00:38.87" lane="2" heatid="18009" points="264" />
                <RESULT resultid="1818" eventid="20" swimtime="00:01:05.98" lane="1" heatid="20022" points="313">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="404" birthdate="2015-01-01" gender="F" lastname="VACOVÁ" firstname="Barbora" license="0">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:44.86" heatid="1003" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:36.20" heatid="7022" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:34.87" heatid="9010" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:44.79" heatid="13008" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:21.74" heatid="19018" lane="2" />
                <ENTRY eventid="21" entrytime="00:03:19.80" heatid="21002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1819" eventid="1" swimtime="00:01:43.06" lane="4" heatid="1003" points="144">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1820" eventid="7" swimtime="00:00:37.23" lane="4" heatid="7022" points="233" />
                <RESULT resultid="1821" eventid="9" swimtime="00:01:35.54" lane="4" heatid="9010" points="206">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1822" eventid="13" swimtime="00:00:44.96" lane="4" heatid="13008" points="159" />
                <RESULT resultid="1823" eventid="19" swimtime="00:01:21.05" lane="2" heatid="19018" points="238">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1824" eventid="21" swimtime="00:03:26.25" lane="3" heatid="21002" points="206">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.26" />
                    <SPLIT distance="100" swimtime="00:01:39.92" />
                    <SPLIT distance="150" swimtime="00:02:43.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="405" birthdate="2017-01-01" gender="M" lastname="VOTRUBEC" firstname="Filip" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:01:12.65" heatid="4001" lane="1" />
                <ENTRY eventid="8" entrytime="00:01:15.00" heatid="8001" lane="1" />
                <ENTRY eventid="16" entrytime="00:02:19.80" heatid="16001" lane="3" />
                <ENTRY eventid="18" entrytime="00:01:22.30" heatid="18001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1825" eventid="4" status="DSQ" swimtime="00:01:12.06" lane="1" heatid="4001" comment="Es erfolgte kein Zielanschlag." />
                <RESULT resultid="1826" eventid="8" swimtime="00:01:23.73" lane="1" heatid="8001" points="13" />
                <RESULT resultid="1827" eventid="16" swimtime="00:02:23.55" lane="3" heatid="16001" points="38" />
                <RESULT resultid="1828" eventid="18" status="DSQ" swimtime="00:01:18.66" lane="1" heatid="18001" comment="Der Sportler startete vor dem Startsignal" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="406" birthdate="2014-01-01" gender="M" lastname="VOTRUBEC" firstname="Tobiás" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:46.82" heatid="4008" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:33.87" heatid="8017" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:28.52" heatid="10006" lane="1" />
                <ENTRY eventid="16" entrytime="00:01:37.88" heatid="16004" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:13.85" heatid="20015" lane="3" />
                <ENTRY eventid="22" entrytime="00:03:36.14" heatid="22002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1829" eventid="4" swimtime="00:00:45.56" lane="4" heatid="4008" points="114" />
                <RESULT resultid="1830" eventid="8" swimtime="00:00:36.16" lane="1" heatid="8017" points="173" />
                <RESULT resultid="1831" eventid="10" swimtime="00:01:32.21" lane="1" heatid="10006" points="152">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1832" eventid="16" swimtime="00:01:35.38" lane="3" heatid="16004" points="130">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1833" eventid="20" swimtime="00:01:15.41" lane="3" heatid="20015" points="210">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1834" eventid="22" swimtime="00:03:15.60" lane="4" heatid="22002" points="176">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:36.26" />
                    <SPLIT distance="150" swimtime="00:02:33.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="407" birthdate="2016-01-01" gender="F" lastname="VOZÁROVÁ" firstname="Alzbeta" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:56.63" heatid="3005" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:42.75" heatid="7012" lane="2" />
                <ENTRY eventid="15" entrytime="00:02:09.46" heatid="15003" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:43.38" heatid="19008" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1835" eventid="3" swimtime="00:00:54.18" lane="3" heatid="3005" points="101" />
                <RESULT resultid="1836" eventid="7" swimtime="00:00:42.72" lane="2" heatid="7012" points="154" />
                <RESULT resultid="1837" eventid="15" swimtime="00:02:00.62" lane="3" heatid="15003" points="94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1838" eventid="19" swimtime="00:01:49.13" lane="4" heatid="19008" points="97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="408" birthdate="2010-01-01" gender="F" lastname="ZELEZNÁ" firstname="Laura" license="0">
              <ENTRIES>
                <ENTRY eventid="29" entrytime="00:01:08.06" heatid="29005" lane="2" />
                <ENTRY eventid="47" entrytime="00:01:12.69" heatid="47006" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:14.81" heatid="33005" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:32.28" heatid="41006" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:05.84" heatid="31011" lane="4" />
                <ENTRY eventid="53" entrytime="00:02:34.63" heatid="53003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1839" eventid="29" swimtime="00:01:13.17" lane="2" heatid="29005" points="403">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1840" eventid="47" swimtime="00:01:15.31" lane="4" heatid="47006" points="387">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1841" eventid="33" swimtime="00:01:15.09" lane="1" heatid="33005" points="426">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1842" eventid="41" swimtime="00:00:32.61" lane="2" heatid="41006" points="417" />
                <RESULT resultid="1843" eventid="31" swimtime="00:01:06.31" lane="4" heatid="31011" points="435">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1844" eventid="53" swimtime="00:02:40.26" lane="1" heatid="53003" points="439">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:02:02.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SSV PCK 90 Schwedt" nation="GER" region="4" code="4738">
          <ATHLETES>
            <ATHLETE athleteid="152" birthdate="2010-01-01" gender="F" lastname="Mau" firstname="Leonie" license="394793" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:25.05" heatid="43012" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:28.13" heatid="41010" lane="2" />
                <ENTRY eventid="25" entrytime="00:00:29.73" heatid="25007" lane="2" />
                <ENTRY eventid="68" entrytime="00:00:25.90" heatid="68001" lane="2" />
                <ENTRY eventid="64" entrytime="00:00:27.72" heatid="64001" lane="2" />
                <ENTRY eventid="56" entrytime="00:00:29.82" heatid="56001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="702" eventid="43" swimtime="00:00:25.90" lane="2" heatid="43012" points="693" />
                <RESULT resultid="703" eventid="41" swimtime="00:00:27.72" lane="2" heatid="41010" points="680" />
                <RESULT resultid="704" eventid="25" swimtime="00:00:29.82" lane="2" heatid="25007" points="607" />
                <RESULT resultid="2351" eventid="56" swimtime="00:00:29.40" lane="2" heatid="56001" points="633" />
                <RESULT resultid="2335" eventid="64" swimtime="00:00:27.76" lane="2" heatid="64001" points="677" />
                <RESULT resultid="2303" eventid="68" swimtime="00:00:25.95" lane="2" heatid="68001" points="689" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="ST Erzgebirge" nation="GER" region="12" code="5134">
          <ATHLETES>
            <ATHLETE athleteid="422" birthdate="2012-01-01" gender="M" lastname="Bochmann" firstname="Noa" license="461952" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:40.33" heatid="4016" lane="4" />
                <ENTRY eventid="6" entrytime="00:01:40.54" heatid="6006" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:34.60" heatid="8016" lane="1" />
                <ENTRY eventid="16" entrytime="00:01:31.17" heatid="16005" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:45.65" heatid="18008" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:14.31" heatid="20015" lane="4" />
                <ENTRY eventid="52" entrytime="00:02:49.15" heatid="52002" lane="1" />
                <ENTRY eventid="36" entrytime="00:03:47.40" heatid="36001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1868" eventid="4" swimtime="00:00:38.47" lane="4" heatid="4016" points="189" />
                <RESULT resultid="1869" eventid="6" status="DSQ" swimtime="00:01:35.50" lane="4" heatid="6006" comment="Beim Zielanschlag hat die Sportlerin mit aufeinandergelegten Händen angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1870" eventid="8" swimtime="00:00:32.47" lane="1" heatid="8016" points="239" />
                <RESULT resultid="1871" eventid="16" swimtime="00:01:31.40" lane="4" heatid="16005" points="147">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1872" eventid="18" swimtime="00:00:44.32" lane="4" heatid="18008" points="178" />
                <RESULT resultid="1873" eventid="20" swimtime="00:01:14.31" lane="4" heatid="20015" points="219">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1874" eventid="52" swimtime="00:02:41.23" lane="1" heatid="52002" points="234">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:58.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1875" eventid="36" swimtime="00:03:14.23" lane="1" heatid="36001" points="160">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                    <SPLIT distance="100" swimtime="00:01:34.03" />
                    <SPLIT distance="150" swimtime="00:02:27.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="423" birthdate="2011-01-01" gender="M" lastname="Fauska" firstname="Franz" license="458123" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:33.38" heatid="44002" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:40.55" heatid="28003" lane="3" />
                <ENTRY eventid="34" entrytime="00:01:25.25" heatid="34002" lane="1" />
                <ENTRY eventid="38" entrytime="00:03:16.00" heatid="38003" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:39.25" heatid="42002" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:28.02" heatid="46004" lane="1" />
                <ENTRY eventid="54" entrytime="00:03:08.79" heatid="54001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1876" eventid="44" swimtime="00:00:32.46" lane="3" heatid="44002" points="239" />
                <RESULT resultid="1877" eventid="28" swimtime="00:00:40.27" lane="3" heatid="28003" points="237" />
                <RESULT resultid="1878" eventid="34" swimtime="00:01:23.07" lane="1" heatid="34002" points="208">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1879" eventid="38" swimtime="00:03:05.52" lane="1" heatid="38003" points="271">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:30.34" />
                    <SPLIT distance="150" swimtime="00:02:18.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1880" eventid="42" swimtime="00:00:39.25" lane="4" heatid="42002" points="170" />
                <RESULT resultid="1881" eventid="46" swimtime="00:01:29.21" lane="1" heatid="46004" points="237">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1882" eventid="54" swimtime="00:03:04.73" lane="3" heatid="54001" points="209">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:01:30.82" />
                    <SPLIT distance="150" swimtime="00:02:21.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="424" birthdate="2013-01-01" gender="F" lastname="Franke" firstname="Jenna" license="497630" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:45.40" heatid="3014" lane="4" />
                <ENTRY eventid="5" entrytime="00:01:43.75" heatid="5008" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:40.47" heatid="7016" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:43.34" heatid="9006" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:47.22" heatid="15007" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:48.39" heatid="17012" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:35.53" heatid="19010" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1883" eventid="3" swimtime="00:00:45.39" lane="4" heatid="3014" points="172" />
                <RESULT resultid="1884" eventid="5" swimtime="00:01:41.42" lane="2" heatid="5008" points="232">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1885" eventid="7" status="DSQ" swimtime="00:00:37.94" lane="4" heatid="7016" comment="Die Sportlerin startete vor dem Startsignal" />
                <RESULT resultid="1886" eventid="9" swimtime="00:01:40.85" lane="4" heatid="9006" points="175">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1887" eventid="15" status="DSQ" swimtime="00:01:44.31" lane="1" heatid="15007" comment="Die Sportlerin hat bei der zweiten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1888" eventid="17" swimtime="00:00:47.76" lane="1" heatid="17012" points="209" />
                <RESULT resultid="1889" eventid="19" swimtime="00:01:30.03" lane="2" heatid="19010" points="173">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="425" birthdate="2011-01-01" gender="M" lastname="Frohs" firstname="Erik" license="480943" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:29.13" heatid="44014" lane="3" />
                <ENTRY eventid="30" entrytime="00:01:15.31" heatid="30003" lane="4" />
                <ENTRY eventid="48" entrytime="00:01:16.43" heatid="48003" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:31.76" heatid="42010" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:34.35" heatid="26007" lane="2" />
                <ENTRY eventid="32" entrytime="00:01:06.36" heatid="32010" lane="1" />
                <ENTRY eventid="54" entrytime="00:02:45.79" heatid="54002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1890" eventid="44" swimtime="00:00:28.70" lane="3" heatid="44014" points="346" />
                <RESULT resultid="1891" eventid="30" swimtime="00:01:11.39" lane="4" heatid="30003" points="299">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1892" eventid="48" swimtime="00:01:20.80" lane="3" heatid="48003" points="214">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1893" eventid="42" swimtime="00:00:30.66" lane="2" heatid="42010" points="356" />
                <RESULT resultid="1894" eventid="26" swimtime="00:00:33.70" lane="2" heatid="26007" points="282" />
                <RESULT resultid="1895" eventid="32" swimtime="00:01:05.52" lane="1" heatid="32010" points="320">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1896" eventid="54" swimtime="00:02:47.82" lane="2" heatid="54002" points="278">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:19.34" />
                    <SPLIT distance="150" swimtime="00:02:09.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="426" birthdate="2017-01-01" gender="F" lastname="Frohs" firstname="Theres" license="511993" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:00.00" heatid="3001" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:51.71" heatid="7005" lane="1" />
                <ENTRY eventid="15" entrytime="00:00:00.00" heatid="15002" lane="1" />
                <ENTRY eventid="19" entrytime="00:02:00.67" heatid="19003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1897" eventid="3" swimtime="00:00:58.54" lane="4" heatid="3001" points="80" />
                <RESULT resultid="1898" eventid="7" swimtime="00:00:52.15" lane="1" heatid="7005" points="85" />
                <RESULT resultid="1899" eventid="15" swimtime="00:02:16.39" lane="1" heatid="15002" points="65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1900" eventid="19" swimtime="00:02:12.45" lane="2" heatid="19003" points="54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="427" birthdate="2009-01-01" gender="M" lastname="Gabler" firstname="Ansgar" license="484404" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:32.64" heatid="44003" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:43.13" heatid="28002" lane="4" />
                <ENTRY eventid="48" entrytime="00:01:26.79" heatid="48001" lane="3" />
                <ENTRY eventid="38" entrytime="00:03:45.91" heatid="38002" lane="1" />
                <ENTRY eventid="26" entrytime="00:00:38.59" heatid="26002" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:38.63" heatid="46001" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:19.13" heatid="32001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1901" eventid="44" swimtime="00:00:32.61" lane="1" heatid="44003" points="236" />
                <RESULT resultid="1902" eventid="28" swimtime="00:00:43.61" lane="4" heatid="28002" points="187" />
                <RESULT resultid="1903" eventid="48" swimtime="00:01:30.25" lane="3" heatid="48001" points="153">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1904" eventid="38" swimtime="00:03:31.01" lane="1" heatid="38002" points="184">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                    <SPLIT distance="100" swimtime="00:01:39.06" />
                    <SPLIT distance="150" swimtime="00:02:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1905" eventid="26" swimtime="00:00:38.67" lane="4" heatid="26002" points="186" />
                <RESULT resultid="1906" eventid="46" swimtime="00:01:37.56" lane="1" heatid="46001" points="181">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1907" eventid="32" swimtime="00:01:22.46" lane="3" heatid="32001" points="160">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="428" birthdate="2013-01-01" gender="M" lastname="Gabler" firstname="Wieland" license="484407" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:46.06" heatid="4008" lane="3" />
                <ENTRY eventid="6" entrytime="00:01:51.25" heatid="6004" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:40.55" heatid="8010" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:45.18" heatid="10002" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:41.69" heatid="16004" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:48.73" heatid="18007" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:36.39" heatid="20006" lane="2" />
                <ENTRY eventid="38" entrytime="00:03:50.86" heatid="38001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1908" eventid="4" swimtime="00:00:44.70" lane="3" heatid="4008" points="121" />
                <RESULT resultid="1909" eventid="6" swimtime="00:01:49.17" lane="4" heatid="6004" points="129">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1910" eventid="8" swimtime="00:00:40.52" lane="3" heatid="8010" points="123" />
                <RESULT resultid="1911" eventid="10" swimtime="00:01:41.44" lane="2" heatid="10002" points="114">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1912" eventid="16" status="DSQ" swimtime="00:01:42.99" lane="4" heatid="16004" comment="Der Sportler hat bei der zweiten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1913" eventid="18" swimtime="00:00:49.48" lane="4" heatid="18007" points="128" />
                <RESULT resultid="1914" eventid="20" swimtime="00:01:31.44" lane="2" heatid="20006" points="117">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1915" eventid="38" swimtime="00:03:55.45" lane="3" heatid="38001" points="132">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.78" />
                    <SPLIT distance="100" swimtime="00:01:52.27" />
                    <SPLIT distance="150" swimtime="00:02:55.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="429" birthdate="2017-01-01" gender="M" lastname="Gimmler" firstname="Hannes" license="505199" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:59.86" heatid="4001" lane="2" />
                <ENTRY eventid="6" entrytime="00:02:15.84" heatid="6007" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:48.12" heatid="8020" lane="1" />
                <ENTRY eventid="18" entrytime="00:01:04.06" heatid="18010" lane="1" />
                <ENTRY eventid="20" entrytime="00:02:02.15" heatid="20001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1916" eventid="4" swimtime="00:00:52.91" lane="2" heatid="4001" points="72" />
                <RESULT resultid="1917" eventid="6" swimtime="00:02:14.93" lane="4" heatid="6007" points="68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1918" eventid="8" swimtime="00:00:46.04" lane="1" heatid="8020" points="83" />
                <RESULT resultid="1919" eventid="18" swimtime="00:01:00.01" lane="1" heatid="18010" points="71" />
                <RESULT resultid="1920" eventid="20" swimtime="00:01:54.36" lane="2" heatid="20001" points="60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="430" birthdate="2012-01-01" gender="M" lastname="Gimmler" firstname="Ruben" license="505198" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:48.21" heatid="4007" lane="1" />
                <ENTRY eventid="6" entrytime="00:01:41.29" heatid="6005" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:34.79" heatid="8015" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:44.63" heatid="18008" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:27.68" heatid="20009" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1921" eventid="4" swimtime="00:00:43.94" lane="1" heatid="4007" points="127" />
                <RESULT resultid="1922" eventid="6" swimtime="00:01:39.50" lane="2" heatid="6005" points="171">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1923" eventid="8" swimtime="00:00:34.66" lane="2" heatid="8015" points="196" />
                <RESULT resultid="1924" eventid="18" swimtime="00:00:44.48" lane="3" heatid="18008" points="176" />
                <RESULT resultid="1925" eventid="20" swimtime="00:01:25.95" lane="3" heatid="20009" points="141">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="431" birthdate="2014-01-01" gender="M" lastname="Gläser" firstname="Julian" license="458122" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:42.39" heatid="4009" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:38.07" heatid="8012" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:37.78" heatid="10004" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:41.97" heatid="14005" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:33.30" heatid="16004" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:27.70" heatid="20009" lane="1" />
                <ENTRY eventid="52" entrytime="00:03:09.47" heatid="52001" lane="3" />
                <ENTRY eventid="36" entrytime="00:03:38.28" heatid="36000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1926" eventid="4" swimtime="00:00:43.69" lane="2" heatid="4009" points="129" />
                <RESULT resultid="1927" eventid="8" swimtime="00:00:37.68" lane="4" heatid="8012" points="153" />
                <RESULT resultid="1928" eventid="10" swimtime="00:01:37.69" lane="1" heatid="10004" points="128">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1929" eventid="14" swimtime="00:00:44.36" lane="3" heatid="14005" points="117" />
                <RESULT resultid="1930" eventid="16" swimtime="00:01:41.62" lane="2" heatid="16004" points="107">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1931" eventid="20" swimtime="00:01:31.18" lane="1" heatid="20009" points="118">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1932" eventid="52" swimtime="00:03:09.90" lane="3" heatid="52001" points="143">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                    <SPLIT distance="100" swimtime="00:01:33.32" />
                    <SPLIT distance="150" swimtime="00:02:24.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1933" eventid="36" status="WDR" swimtime="00:00:00.00" lane="0" heatid="36000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="432" birthdate="2010-01-01" gender="M" lastname="Gläser" firstname="Simon" license="461951" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:30.91" heatid="44004" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:39.96" heatid="28003" lane="2" />
                <ENTRY eventid="34" entrytime="00:01:19.84" heatid="34003" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:35.97" heatid="42003" lane="3" />
                <ENTRY eventid="46" entrytime="00:01:26.85" heatid="46001" lane="2" />
                <ENTRY eventid="32" entrytime="00:01:12.44" heatid="32003" lane="4" />
                <ENTRY eventid="54" entrytime="00:03:00.23" heatid="54002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1934" eventid="44" swimtime="00:00:30.98" lane="4" heatid="44004" points="275" />
                <RESULT resultid="1935" eventid="28" swimtime="00:00:37.58" lane="2" heatid="28003" points="292" />
                <RESULT resultid="1936" eventid="34" swimtime="00:01:20.44" lane="2" heatid="34003" points="229">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1937" eventid="42" swimtime="00:00:36.66" lane="3" heatid="42003" points="208" />
                <RESULT resultid="1938" eventid="46" swimtime="00:01:27.22" lane="2" heatid="46001" points="254">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1939" eventid="32" swimtime="00:01:14.29" lane="4" heatid="32003" points="219">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1940" eventid="54" swimtime="00:03:04.08" lane="4" heatid="54002" points="211">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:26.44" />
                    <SPLIT distance="150" swimtime="00:02:18.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="433" birthdate="2017-01-01" gender="F" lastname="Glöckner" firstname="Tia" license="511997" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:01:00.06" heatid="3002" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:53.62" heatid="7005" lane="4" />
                <ENTRY eventid="9" entrytime="00:00:00.00" heatid="9001" lane="3" />
                <ENTRY eventid="15" entrytime="00:00:00.00" heatid="15001" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:00.00" heatid="17001" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:50.69" heatid="19004" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1941" eventid="3" swimtime="00:00:53.71" lane="2" heatid="3002" points="103" />
                <RESULT resultid="1942" eventid="7" swimtime="00:00:56.10" lane="4" heatid="7005" points="68" />
                <RESULT resultid="1943" eventid="9" swimtime="00:02:32.93" lane="3" heatid="9001" points="50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1944" eventid="15" swimtime="00:02:11.12" lane="2" heatid="15001" points="73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1945" eventid="17" swimtime="00:01:11.19" lane="1" heatid="17001" points="63" />
                <RESULT resultid="1946" eventid="19" swimtime="00:02:12.12" lane="2" heatid="19004" points="55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="434" birthdate="2010-01-01" gender="F" lastname="Göhler" firstname="Lucy" license="402479" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:31.41" heatid="43007" lane="4" />
                <ENTRY eventid="47" entrytime="00:01:20.07" heatid="47002" lane="2" />
                <ENTRY eventid="51" entrytime="00:02:34.03" heatid="51002" lane="1" />
                <ENTRY eventid="25" entrytime="00:00:34.91" heatid="25004" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:09.05" heatid="31007" lane="3" />
                <ENTRY eventid="53" entrytime="00:02:53.20" heatid="53002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1947" eventid="43" swimtime="00:00:31.89" lane="4" heatid="43007" points="371" />
                <RESULT resultid="1948" eventid="47" swimtime="00:01:18.38" lane="2" heatid="47002" points="343">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1949" eventid="51" swimtime="00:02:32.13" lane="1" heatid="51002" points="381">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:01:52.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1950" eventid="25" swimtime="00:00:35.82" lane="1" heatid="25004" points="350" />
                <RESULT resultid="1951" eventid="31" swimtime="00:01:09.83" lane="3" heatid="31007" points="372">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1952" eventid="53" swimtime="00:02:53.64" lane="1" heatid="53002" points="345">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:23.49" />
                    <SPLIT distance="150" swimtime="00:02:14.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="435" birthdate="2012-01-01" gender="M" lastname="Gottschalk" firstname="Karl" license="461957" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:46.15" heatid="4008" lane="1" />
                <ENTRY eventid="6" entrytime="00:01:41.57" heatid="6005" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:35.66" heatid="8014" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:38.38" heatid="10003" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:46.16" heatid="14004" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:44.10" heatid="18009" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:23.66" heatid="20011" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1953" eventid="4" swimtime="00:00:45.73" lane="1" heatid="4008" points="113" />
                <RESULT resultid="1954" eventid="6" swimtime="00:01:36.26" lane="3" heatid="6005" points="189">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1955" eventid="8" swimtime="00:00:34.86" lane="3" heatid="8014" points="193" />
                <RESULT resultid="1956" eventid="10" swimtime="00:01:32.82" lane="2" heatid="10003" points="149">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1957" eventid="14" swimtime="00:00:44.76" lane="1" heatid="14004" points="114" />
                <RESULT resultid="1958" eventid="18" swimtime="00:00:43.93" lane="1" heatid="18009" points="183" />
                <RESULT resultid="1959" eventid="20" swimtime="00:01:22.96" lane="1" heatid="20011" points="157">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="437" birthdate="2013-01-01" gender="F" lastname="Günther" firstname="Zoe-Marie" license="497632" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:48.84" heatid="3010" lane="1" />
                <ENTRY eventid="5" entrytime="00:01:53.65" heatid="5005" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:42.43" heatid="7013" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:50.53" heatid="13004" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:50.81" heatid="17010" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:37.65" heatid="19009" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1963" eventid="3" swimtime="00:00:47.73" lane="1" heatid="3010" points="148" />
                <RESULT resultid="1964" eventid="5" swimtime="00:01:57.11" lane="3" heatid="5005" points="150">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1965" eventid="7" swimtime="00:00:43.25" lane="3" heatid="7013" points="149" />
                <RESULT resultid="1966" eventid="13" swimtime="00:00:52.57" lane="1" heatid="13004" points="99" />
                <RESULT resultid="1967" eventid="17" swimtime="00:00:54.23" lane="2" heatid="17010" points="143" />
                <RESULT resultid="1968" eventid="19" swimtime="00:01:36.58" lane="2" heatid="19009" points="140">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="438" birthdate="2017-01-01" gender="F" lastname="Haufe-Reichel" firstname="Leni" license="511996" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:01:00.18" heatid="3002" lane="3" />
                <ENTRY eventid="5" entrytime="00:02:17.93" heatid="5002" lane="2" />
                <ENTRY eventid="7" entrytime="00:01:01.05" heatid="7001" lane="2" />
                <ENTRY eventid="15" entrytime="00:02:08.90" heatid="15003" lane="2" />
                <ENTRY eventid="17" entrytime="00:01:02.85" heatid="17004" lane="1" />
                <ENTRY eventid="19" entrytime="00:00:00.00" heatid="19001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1969" eventid="3" swimtime="00:00:55.49" lane="3" heatid="3002" points="94" />
                <RESULT resultid="1970" eventid="5" swimtime="00:02:16.36" lane="2" heatid="5002" points="95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1971" eventid="7" swimtime="00:00:55.06" lane="2" heatid="7001" points="72" />
                <RESULT resultid="1972" eventid="15" swimtime="00:02:04.02" lane="2" heatid="15003" points="86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1973" eventid="17" swimtime="00:01:02.60" lane="1" heatid="17004" points="93" />
                <RESULT resultid="1974" eventid="19" swimtime="00:02:05.18" lane="1" heatid="19001" points="64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="439" birthdate="2011-01-01" gender="F" lastname="Hiemann" firstname="Elisa" license="461993" nation="GER">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:39.85" heatid="27007" lane="3" />
                <ENTRY eventid="29" entrytime="00:01:19.41" heatid="29004" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:21.33" heatid="33007" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:33.53" heatid="41009" lane="3" />
                <ENTRY eventid="45" entrytime="00:01:26.95" heatid="45005" lane="3" />
                <ENTRY eventid="53" entrytime="00:03:00.93" heatid="53001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1975" eventid="27" swimtime="00:00:38.52" lane="3" heatid="27007" points="399" />
                <RESULT resultid="1976" eventid="29" swimtime="00:01:18.16" lane="2" heatid="29004" points="330">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1977" eventid="33" swimtime="00:01:19.78" lane="4" heatid="33007" points="355">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1978" eventid="41" swimtime="00:00:33.56" lane="3" heatid="41009" points="383" />
                <RESULT resultid="1979" eventid="45" swimtime="00:01:26.92" lane="3" heatid="45005" points="369">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1980" eventid="53" swimtime="00:02:52.38" lane="1" heatid="53001" points="353">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:09.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="440" birthdate="2016-01-01" gender="M" lastname="Hiemann" firstname="Erik" license="490703" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:46.64" heatid="6008" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:46.82" heatid="8005" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:51.45" heatid="10009" lane="4" />
                <ENTRY eventid="14" entrytime="00:00:55.99" heatid="14002" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:47.67" heatid="18011" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:49.99" heatid="20003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1981" eventid="6" swimtime="00:01:41.31" lane="2" heatid="6008" points="162">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1982" eventid="8" swimtime="00:00:42.74" lane="4" heatid="8005" points="104" />
                <RESULT resultid="1983" eventid="10" swimtime="00:01:51.35" lane="4" heatid="10009" points="86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1984" eventid="14" swimtime="00:01:02.16" lane="3" heatid="14002" points="42" />
                <RESULT resultid="1985" eventid="18" swimtime="00:00:48.21" lane="2" heatid="18011" points="138" />
                <RESULT resultid="1986" eventid="20" swimtime="00:01:40.10" lane="1" heatid="20003" points="89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="441" birthdate="2014-01-01" gender="F" lastname="Hübler" firstname="Laureen" license="497633" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:58.09" heatid="3004" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:50.49" heatid="7006" lane="2" />
                <ENTRY eventid="17" entrytime="00:01:02.11" heatid="17004" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1987" eventid="3" swimtime="00:00:53.35" lane="2" heatid="3004" points="106" />
                <RESULT resultid="1988" eventid="7" swimtime="00:00:45.46" lane="2" heatid="7006" points="128" />
                <RESULT resultid="1989" eventid="17" swimtime="00:00:57.18" lane="3" heatid="17004" points="122" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="442" birthdate="2011-01-01" gender="F" lastname="Kaden" firstname="Nele" license="466489" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:36.88" heatid="43000" lane="0" />
                <ENTRY eventid="47" entrytime="00:01:38.99" heatid="47000" lane="0" />
                <ENTRY eventid="41" entrytime="00:00:43.89" heatid="41000" lane="0" />
                <ENTRY eventid="25" entrytime="00:00:43.80" heatid="25000" lane="0" />
                <ENTRY eventid="31" entrytime="00:01:26.52" heatid="31000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1990" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
                <RESULT resultid="1991" eventid="47" status="WDR" swimtime="00:00:00.00" lane="0" heatid="47000" />
                <RESULT resultid="1992" eventid="41" status="WDR" swimtime="00:00:00.00" lane="0" heatid="41000" />
                <RESULT resultid="1993" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
                <RESULT resultid="1994" eventid="31" status="WDR" swimtime="00:00:00.00" lane="0" heatid="31000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="443" birthdate="2002-01-01" gender="F" lastname="Katsala" firstname="Mariia" license="458276" nation="UKR">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:31.66" heatid="43000" lane="0" />
                <ENTRY eventid="47" entrytime="00:01:09.20" heatid="47000" lane="0" />
                <ENTRY eventid="25" entrytime="00:00:33.98" heatid="25000" lane="0" />
                <ENTRY eventid="31" entrytime="00:01:05.56" heatid="31000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1995" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
                <RESULT resultid="1996" eventid="47" status="WDR" swimtime="00:00:00.00" lane="0" heatid="47000" />
                <RESULT resultid="1997" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
                <RESULT resultid="1998" eventid="31" status="WDR" swimtime="00:00:00.00" lane="0" heatid="31000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="444" birthdate="2014-01-01" gender="M" lastname="Kirsche" firstname="Linus" license="500601" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:48.96" heatid="4006" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:53.70" heatid="8002" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:00.00" heatid="14001" lane="1" />
                <ENTRY eventid="16" entrytime="00:02:03.42" heatid="16001" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:55.84" heatid="20002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1999" eventid="4" swimtime="00:00:48.25" lane="2" heatid="4006" points="96" />
                <RESULT resultid="2000" eventid="8" swimtime="00:00:47.08" lane="2" heatid="8002" points="78" />
                <RESULT resultid="2001" eventid="14" swimtime="00:00:59.65" lane="1" heatid="14001" points="48" />
                <RESULT resultid="2002" eventid="16" swimtime="00:01:49.13" lane="2" heatid="16001" points="86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2003" eventid="20" swimtime="00:01:47.18" lane="1" heatid="20002" points="73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="445" birthdate="2013-01-01" gender="F" lastname="Klaus" firstname="Emma" license="461960" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.74" heatid="3014" lane="3" />
                <ENTRY eventid="5" entrytime="00:01:43.41" heatid="5009" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:36.63" heatid="7021" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:35.32" heatid="9009" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:46.23" heatid="13007" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:46.04" heatid="17014" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:27.04" heatid="19014" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2004" eventid="3" swimtime="00:00:44.47" lane="3" heatid="3014" points="183" />
                <RESULT resultid="2005" eventid="5" swimtime="00:01:49.32" lane="3" heatid="5009" points="185">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2006" eventid="7" swimtime="00:00:36.35" lane="4" heatid="7021" points="251" />
                <RESULT resultid="2007" eventid="9" swimtime="00:01:34.23" lane="2" heatid="9009" points="215">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2008" eventid="13" swimtime="00:00:46.18" lane="4" heatid="13007" points="147" />
                <RESULT resultid="2009" eventid="17" swimtime="00:00:48.01" lane="2" heatid="17014" points="206" />
                <RESULT resultid="2010" eventid="19" swimtime="00:01:27.24" lane="3" heatid="19014" points="191">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="446" birthdate="2013-01-01" gender="M" lastname="Konrad" firstname="Christian" license="461953" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:35.88" heatid="2002" lane="1" />
                <ENTRY eventid="6" entrytime="00:01:31.84" heatid="6011" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:33.99" heatid="8017" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:26.00" heatid="10007" lane="4" />
                <ENTRY eventid="14" entrytime="00:00:38.41" heatid="14006" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:40.77" heatid="18014" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:17.77" heatid="20013" lane="4" />
                <ENTRY eventid="38" entrytime="00:03:23.65" heatid="38003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2011" eventid="2" swimtime="00:01:37.44" lane="1" heatid="2002" points="117">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2012" eventid="6" swimtime="00:01:30.76" lane="3" heatid="6011" points="225">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2013" eventid="8" swimtime="00:00:34.11" lane="4" heatid="8017" points="206" />
                <RESULT resultid="2014" eventid="10" swimtime="00:01:25.12" lane="4" heatid="10007" points="194">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2015" eventid="14" swimtime="00:00:40.82" lane="1" heatid="14006" points="151" />
                <RESULT resultid="2016" eventid="18" swimtime="00:00:41.88" lane="1" heatid="18014" points="211" />
                <RESULT resultid="2017" eventid="20" swimtime="00:01:21.40" lane="4" heatid="20013" points="167">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2018" eventid="38" swimtime="00:03:20.04" lane="4" heatid="38003" points="216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                    <SPLIT distance="100" swimtime="00:01:37.70" />
                    <SPLIT distance="150" swimtime="00:02:30.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="447" birthdate="2008-01-01" gender="M" lastname="Kulai" firstname="Vasyl" license="429668" nation="UKR">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:37.28" heatid="28004" lane="2" />
                <ENTRY eventid="48" entrytime="00:01:21.56" heatid="48002" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:20.86" heatid="34003" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:35.40" heatid="26003" lane="3" />
                <ENTRY eventid="46" entrytime="00:01:22.39" heatid="46002" lane="3" />
                <ENTRY eventid="54" entrytime="00:02:56.42" heatid="54002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2019" eventid="28" swimtime="00:00:36.23" lane="2" heatid="28004" points="326" />
                <RESULT resultid="2020" eventid="48" swimtime="00:01:20.65" lane="1" heatid="48002" points="215">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2021" eventid="34" swimtime="00:01:15.59" lane="4" heatid="34003" points="277">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2022" eventid="26" swimtime="00:00:36.51" lane="3" heatid="26003" points="222" />
                <RESULT resultid="2023" eventid="46" swimtime="00:01:22.55" lane="3" heatid="46002" points="300">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2024" eventid="54" swimtime="00:02:52.25" lane="1" heatid="54002" points="257">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:21.80" />
                    <SPLIT distance="150" swimtime="00:02:08.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="448" birthdate="2015-01-01" gender="F" lastname="Kunze" firstname="Ella" license="490707" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:49.30" heatid="3010" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:44.22" heatid="7011" lane="4" />
                <ENTRY eventid="9" entrytime="00:00:00.00" heatid="9001" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:56.23" heatid="13002" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:50.52" heatid="15006" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:40.08" heatid="19009" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2025" eventid="3" swimtime="00:00:48.09" lane="4" heatid="3010" points="144" />
                <RESULT resultid="2026" eventid="7" swimtime="00:00:44.34" lane="4" heatid="7011" points="138" />
                <RESULT resultid="2027" eventid="9" swimtime="00:01:49.18" lane="1" heatid="9001" points="138">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2028" eventid="13" swimtime="00:00:51.82" lane="2" heatid="13002" points="104" />
                <RESULT resultid="2029" eventid="15" swimtime="00:01:47.22" lane="1" heatid="15006" points="134">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2030" eventid="19" swimtime="00:01:41.09" lane="4" heatid="19009" points="122">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="449" birthdate="2012-01-01" gender="F" lastname="Langer" firstname="Mia" license="461959" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:37.69" heatid="43001" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:46.66" heatid="27002" lane="1" />
                <ENTRY eventid="47" entrytime="00:01:51.42" heatid="47004" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:38.16" heatid="33001" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:45.34" heatid="41001" lane="1" />
                <ENTRY eventid="25" entrytime="00:00:44.79" heatid="25001" lane="3" />
                <ENTRY eventid="45" entrytime="00:01:47.80" heatid="45001" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:26.05" heatid="31001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2031" eventid="43" swimtime="00:00:36.04" lane="2" heatid="43001" points="257" />
                <RESULT resultid="2032" eventid="27" swimtime="00:00:44.83" lane="1" heatid="27002" points="253" />
                <RESULT resultid="2033" eventid="47" swimtime="00:01:37.47" lane="4" heatid="47004" points="178">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2034" eventid="33" swimtime="00:01:37.40" lane="2" heatid="33001" points="195">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2035" eventid="41" swimtime="00:00:41.37" lane="1" heatid="41001" points="204" />
                <RESULT resultid="2036" eventid="25" swimtime="00:00:44.07" lane="3" heatid="25001" points="188" />
                <RESULT resultid="2037" eventid="45" swimtime="00:01:45.13" lane="3" heatid="45001" points="208">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2038" eventid="31" swimtime="00:01:27.42" lane="2" heatid="31001" points="189">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="450" birthdate="2013-01-01" gender="M" lastname="Langer" firstname="Paul" license="480942" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:44.43" heatid="4008" lane="2" />
                <ENTRY eventid="6" entrytime="00:01:37.60" heatid="6011" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:35.16" heatid="8015" lane="4" />
                <ENTRY eventid="14" entrytime="00:00:46.33" heatid="14004" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:45.31" heatid="18008" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:23.38" heatid="20011" lane="3" />
                <ENTRY eventid="38" entrytime="00:03:50.79" heatid="38001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2039" eventid="4" swimtime="00:00:43.25" lane="2" heatid="4008" points="133" />
                <RESULT resultid="2040" eventid="6" swimtime="00:01:33.58" lane="1" heatid="6011" points="206">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2041" eventid="8" swimtime="00:00:34.81" lane="4" heatid="8015" points="194" />
                <RESULT resultid="2042" eventid="14" swimtime="00:00:38.36" lane="4" heatid="14004" points="182" />
                <RESULT resultid="2043" eventid="18" swimtime="00:00:43.61" lane="1" heatid="18008" points="187" />
                <RESULT resultid="2044" eventid="20" swimtime="00:01:19.85" lane="3" heatid="20011" points="177">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2045" eventid="38" swimtime="00:03:24.74" lane="2" heatid="38001" points="202">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.50" />
                    <SPLIT distance="100" swimtime="00:01:40.00" />
                    <SPLIT distance="150" swimtime="00:02:33.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="451" birthdate="2013-01-01" gender="M" lastname="Lehmann" firstname="Jay" license="461955" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:49.00" heatid="2001" lane="1" />
                <ENTRY eventid="4" entrytime="00:00:46.90" heatid="4007" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:40.55" heatid="8010" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:40.77" heatid="10003" lane="4" />
                <ENTRY eventid="14" entrytime="00:00:46.03" heatid="14004" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:30.27" heatid="20008" lane="3" />
                <ENTRY eventid="52" entrytime="00:03:14.54" heatid="52001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2046" eventid="2" swimtime="00:01:52.21" lane="1" heatid="2001" points="77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2047" eventid="4" swimtime="00:00:46.59" lane="2" heatid="4007" points="106" />
                <RESULT resultid="2048" eventid="8" swimtime="00:00:39.93" lane="1" heatid="8010" points="128" />
                <RESULT resultid="2049" eventid="10" swimtime="00:01:41.97" lane="4" heatid="10003" points="112">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2050" eventid="14" swimtime="00:00:51.02" lane="3" heatid="14004" points="77" />
                <RESULT resultid="2051" eventid="20" swimtime="00:01:30.20" lane="3" heatid="20008" points="122">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2052" eventid="52" swimtime="00:03:08.59" lane="1" heatid="52001" points="146">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:30.56" />
                    <SPLIT distance="150" swimtime="00:02:18.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="452" birthdate="2010-01-01" gender="F" lastname="Lorenz" firstname="Milena" license="417871" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:35.23" heatid="43003" lane="4" />
                <ENTRY eventid="29" entrytime="00:01:32.81" heatid="29001" lane="2" />
                <ENTRY eventid="47" entrytime="00:01:37.51" heatid="47001" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:39.22" heatid="41003" lane="1" />
                <ENTRY eventid="25" entrytime="00:00:42.53" heatid="25002" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:20.56" heatid="31002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2053" eventid="43" swimtime="00:00:34.85" lane="4" heatid="43003" points="284" />
                <RESULT resultid="2054" eventid="29" swimtime="00:01:35.97" lane="2" heatid="29001" points="178">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2055" eventid="47" swimtime="00:01:41.11" lane="3" heatid="47001" points="159">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2056" eventid="41" swimtime="00:00:39.96" lane="1" heatid="41003" points="227" />
                <RESULT resultid="2057" eventid="25" swimtime="00:00:44.78" lane="4" heatid="25002" points="179" />
                <RESULT resultid="2058" eventid="31" swimtime="00:01:22.13" lane="3" heatid="31002" points="229">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="453" birthdate="2016-01-01" gender="F" lastname="Meyer" firstname="Lilly" license="490705" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:00:00.00" heatid="5001" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:54.86" heatid="7004" lane="1" />
                <ENTRY eventid="17" entrytime="00:01:00.99" heatid="17005" lane="1" />
                <ENTRY eventid="19" entrytime="00:00:00.00" heatid="19001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2059" eventid="5" swimtime="00:02:13.07" lane="3" heatid="5001" points="102">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2060" eventid="7" swimtime="00:00:49.63" lane="1" heatid="7004" points="98" />
                <RESULT resultid="2061" eventid="17" swimtime="00:01:02.44" lane="1" heatid="17005" points="93" />
                <RESULT resultid="2062" eventid="19" swimtime="00:02:00.12" lane="2" heatid="19001" points="73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="454" birthdate="2013-01-01" gender="M" lastname="Meyer" firstname="Sammy" license="458126" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:37.80" heatid="4015" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:33.03" heatid="8018" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:29.40" heatid="10006" lane="4" />
                <ENTRY eventid="14" entrytime="00:00:39.08" heatid="14006" lane="4" />
                <ENTRY eventid="16" entrytime="00:01:25.57" heatid="16010" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:14.24" heatid="20015" lane="1" />
                <ENTRY eventid="22" entrytime="00:03:17.85" heatid="22002" lane="2" />
                <ENTRY eventid="52" entrytime="00:02:46.78" heatid="52002" lane="3" />
                <ENTRY eventid="36" entrytime="00:03:02.74" heatid="36001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2063" eventid="4" swimtime="00:00:35.43" lane="3" heatid="4015" points="243" />
                <RESULT resultid="2064" eventid="8" swimtime="00:00:30.84" lane="3" heatid="8018" points="279" />
                <RESULT resultid="2065" eventid="10" swimtime="00:01:23.13" lane="4" heatid="10006" points="208">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2066" eventid="14" swimtime="00:00:36.87" lane="4" heatid="14006" points="205" />
                <RESULT resultid="2067" eventid="16" swimtime="00:01:23.23" lane="3" heatid="16010" points="195">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2068" eventid="20" swimtime="00:01:12.67" lane="1" heatid="20015" points="234">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2069" eventid="22" swimtime="00:03:05.49" lane="2" heatid="22002" points="206">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:30.31" />
                    <SPLIT distance="150" swimtime="00:02:25.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2070" eventid="52" swimtime="00:02:36.34" lane="3" heatid="52002" points="256">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:15.67" />
                    <SPLIT distance="150" swimtime="00:01:57.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2071" eventid="36" swimtime="00:02:59.75" lane="3" heatid="36001" points="202">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                    <SPLIT distance="100" swimtime="00:01:28.64" />
                    <SPLIT distance="150" swimtime="00:02:15.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="455" birthdate="2013-01-01" gender="F" lastname="Mildner" firstname="Donna" license="480945" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:43.25" heatid="1005" lane="4" />
                <ENTRY eventid="3" entrytime="00:00:43.17" heatid="3016" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:36.84" heatid="7020" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:36.65" heatid="9008" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:43.30" heatid="13009" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:38.05" heatid="15010" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:26.56" heatid="19014" lane="2" />
                <ENTRY eventid="51" entrytime="00:03:06.44" heatid="51000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2072" eventid="1" status="DNS" swimtime="00:00:00.00" lane="4" heatid="1005" />
                <RESULT resultid="2073" eventid="3" status="DNS" swimtime="00:00:00.00" lane="1" heatid="3016" />
                <RESULT resultid="2074" eventid="7" status="DNS" swimtime="00:00:00.00" lane="2" heatid="7020" />
                <RESULT resultid="2075" eventid="9" status="DNS" swimtime="00:00:00.00" lane="3" heatid="9008" />
                <RESULT resultid="2076" eventid="13" status="DNS" swimtime="00:00:00.00" lane="1" heatid="13009" />
                <RESULT resultid="2077" eventid="15" status="DNS" swimtime="00:00:00.00" lane="3" heatid="15010" />
                <RESULT resultid="2078" eventid="19" status="DNS" swimtime="00:00:00.00" lane="2" heatid="19014" />
                <RESULT resultid="2079" eventid="51" status="WDR" swimtime="00:00:00.00" lane="0" heatid="51000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="456" birthdate="2015-01-01" gender="F" lastname="Morgenstern" firstname="Elena" license="471532" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:47.61" heatid="3000" lane="0" />
                <ENTRY eventid="5" entrytime="00:01:45.14" heatid="5000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:40.41" heatid="7000" lane="0" />
                <ENTRY eventid="9" entrytime="00:01:53.21" heatid="9000" lane="0" />
                <ENTRY eventid="17" entrytime="00:00:47.88" heatid="17000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:45.99" heatid="19000" lane="0" />
                <ENTRY eventid="37" entrytime="00:00:00.00" heatid="37000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2080" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="2081" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="2082" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="2083" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
                <RESULT resultid="2084" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
                <RESULT resultid="2085" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
                <RESULT resultid="2086" eventid="37" status="WDR" swimtime="00:00:00.00" lane="0" heatid="37000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="457" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Annica" license="429663" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:31.09" heatid="43011" lane="1" />
                <ENTRY eventid="29" entrytime="00:01:22.99" heatid="29004" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:22.35" heatid="33004" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:34.15" heatid="41009" lane="1" />
                <ENTRY eventid="25" entrytime="00:00:37.68" heatid="25006" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:09.83" heatid="31010" lane="1" />
                <ENTRY eventid="53" entrytime="00:03:03.07" heatid="53001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2087" eventid="43" swimtime="00:00:31.28" lane="1" heatid="43011" points="393" />
                <RESULT resultid="2088" eventid="29" swimtime="00:01:21.62" lane="3" heatid="29004" points="290">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2089" eventid="33" swimtime="00:01:21.18" lane="1" heatid="33004" points="337">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2090" eventid="41" swimtime="00:00:34.74" lane="1" heatid="41009" points="345" />
                <RESULT resultid="2091" eventid="25" swimtime="00:00:38.02" lane="4" heatid="25006" points="292" />
                <RESULT resultid="2092" eventid="31" swimtime="00:01:09.00" lane="1" heatid="31010" points="386">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2093" eventid="53" swimtime="00:02:56.56" lane="4" heatid="53001" points="328">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:21.93" />
                    <SPLIT distance="150" swimtime="00:02:13.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="458" birthdate="2012-01-01" gender="F" lastname="Müller" firstname="Frida" license="461992" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:33.44" heatid="43005" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:45.08" heatid="27002" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:26.46" heatid="33006" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:37.49" heatid="41008" lane="4" />
                <ENTRY eventid="45" entrytime="00:01:35.74" heatid="45004" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:15.97" heatid="31004" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2094" eventid="43" swimtime="00:00:32.99" lane="4" heatid="43005" points="335" />
                <RESULT resultid="2095" eventid="27" swimtime="00:00:45.94" lane="3" heatid="27002" points="235" />
                <RESULT resultid="2096" eventid="33" swimtime="00:01:25.89" lane="4" heatid="33006" points="284">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2097" eventid="41" swimtime="00:00:36.48" lane="4" heatid="41008" points="298" />
                <RESULT resultid="2098" eventid="45" swimtime="00:01:38.93" lane="1" heatid="45004" points="250">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2099" eventid="31" swimtime="00:01:15.02" lane="3" heatid="31004" points="300">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="459" birthdate="2009-01-01" gender="M" lastname="Neubert" firstname="Domenic" license="429667" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.98" heatid="44002" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:31.45" heatid="42001" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:24.51" heatid="46004" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:04.85" heatid="32001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2100" eventid="44" swimtime="00:00:27.62" lane="4" heatid="44002" points="388" />
                <RESULT resultid="2102" eventid="42" status="DSQ" swimtime="00:00:30.95" lane="4" heatid="42001" comment="Der Sportler führte mit den Beinen wechselseitig Bewegungen aus." />
                <RESULT resultid="2103" eventid="46" swimtime="00:01:25.47" lane="4" heatid="46004" points="270">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2104" eventid="32" swimtime="00:01:08.47" lane="4" heatid="32001" points="280">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="460" birthdate="2016-01-01" gender="F" lastname="Neubert" firstname="Lissi" license="490704" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:01:03.69" heatid="3002" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:49.52" heatid="7007" lane="2" />
                <ENTRY eventid="9" entrytime="00:00:00.00" heatid="9001" lane="2" />
                <ENTRY eventid="13" entrytime="00:01:08.28" heatid="13001" lane="3" />
                <ENTRY eventid="15" entrytime="00:02:27.18" heatid="15003" lane="1" />
                <ENTRY eventid="19" entrytime="00:02:03.39" heatid="19002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2105" eventid="3" swimtime="00:00:58.91" lane="4" heatid="3002" points="78" />
                <RESULT resultid="2106" eventid="7" swimtime="00:00:46.63" lane="2" heatid="7007" points="118" />
                <RESULT resultid="2107" eventid="9" swimtime="00:02:05.16" lane="2" heatid="9001" points="92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2108" eventid="13" swimtime="00:01:01.01" lane="3" heatid="13001" points="63" />
                <RESULT resultid="2109" eventid="15" swimtime="00:02:19.07" lane="1" heatid="15003" points="61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2110" eventid="19" swimtime="00:01:54.77" lane="2" heatid="19002" points="83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="461" birthdate="2013-01-01" gender="M" lastname="Nordheim" firstname="Matteo" license="461956" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:48.12" heatid="4007" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:40.40" heatid="8010" lane="2" />
                <ENTRY eventid="10" entrytime="00:00:00.00" heatid="10001" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:47.89" heatid="14003" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:41.84" heatid="16003" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:29.40" heatid="20008" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2111" eventid="4" status="DNS" swimtime="00:00:00.00" lane="3" heatid="4007" />
                <RESULT resultid="2112" eventid="8" status="DNS" swimtime="00:00:00.00" lane="2" heatid="8010" />
                <RESULT resultid="2113" eventid="10" status="DNS" swimtime="00:00:00.00" lane="1" heatid="10001" />
                <RESULT resultid="2114" eventid="14" status="DNS" swimtime="00:00:00.00" lane="2" heatid="14003" />
                <RESULT resultid="2115" eventid="16" status="DNS" swimtime="00:00:00.00" lane="2" heatid="16003" />
                <RESULT resultid="2116" eventid="20" status="DNS" swimtime="00:00:00.00" lane="2" heatid="20008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="462" birthdate="2016-01-01" gender="F" lastname="Oestreich" firstname="Leonie" license="490897" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.60" heatid="3020" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:40.14" heatid="7016" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:45.35" heatid="9004" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:39.13" heatid="15016" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:50.45" heatid="17017" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:31.66" heatid="19013" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2117" eventid="3" swimtime="00:00:45.17" lane="1" heatid="3020" points="174" />
                <RESULT resultid="2118" eventid="7" swimtime="00:00:39.96" lane="3" heatid="7016" points="188" />
                <RESULT resultid="2119" eventid="9" swimtime="00:01:40.35" lane="2" heatid="9004" points="178">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2120" eventid="15" swimtime="00:01:42.31" lane="3" heatid="15016" points="154">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2121" eventid="17" swimtime="00:00:51.74" lane="1" heatid="17017" points="164" />
                <RESULT resultid="2122" eventid="19" swimtime="00:01:34.09" lane="1" heatid="19013" points="152">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="463" birthdate="2013-01-01" gender="F" lastname="Oestreich" firstname="Sophia" license="458275" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:40.43" heatid="3018" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:36.15" heatid="7022" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:38.66" heatid="9006" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:28.76" heatid="15013" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:24.03" heatid="19016" lane="4" />
                <ENTRY eventid="51" entrytime="00:03:08.00" heatid="51001" lane="1" />
                <ENTRY eventid="35" entrytime="00:03:28.24" heatid="35001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2123" eventid="3" swimtime="00:00:40.00" lane="1" heatid="3018" points="251" />
                <RESULT resultid="2124" eventid="7" swimtime="00:00:34.34" lane="3" heatid="7022" points="297" />
                <RESULT resultid="2125" eventid="9" swimtime="00:01:34.45" lane="2" heatid="9006" points="214">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2126" eventid="15" swimtime="00:01:34.28" lane="2" heatid="15013" points="197">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2127" eventid="19" swimtime="00:01:22.84" lane="4" heatid="19016" points="223">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2128" eventid="51" swimtime="00:03:01.15" lane="1" heatid="51001" points="225">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.72" />
                    <SPLIT distance="150" swimtime="00:02:13.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2129" eventid="35" status="DSQ" swimtime="00:03:16.62" lane="1" heatid="35001" comment="Bei der sechsten Wende hat die Sportlerin die Wand verlassen, bevor die Rückenlage eingenommen war.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                    <SPLIT distance="100" swimtime="00:01:33.80" />
                    <SPLIT distance="150" swimtime="00:02:24.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="464" birthdate="2014-01-01" gender="F" lastname="Popp" firstname="Hanna" license="511995" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:00.00" heatid="3001" lane="1" />
                <ENTRY eventid="5" entrytime="00:01:56.55" heatid="5004" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:00.00" heatid="7001" lane="1" />
                <ENTRY eventid="15" entrytime="00:00:00.00" heatid="15002" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:52.17" heatid="17009" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2130" eventid="3" swimtime="00:00:53.25" lane="1" heatid="3001" points="106" />
                <RESULT resultid="2131" eventid="5" swimtime="00:01:55.29" lane="2" heatid="5004" points="158">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2132" eventid="7" swimtime="00:00:53.21" lane="1" heatid="7001" points="80" />
                <RESULT resultid="2133" eventid="15" swimtime="00:02:05.58" lane="2" heatid="15002" points="83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2134" eventid="17" swimtime="00:00:56.13" lane="2" heatid="17009" points="129" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="465" birthdate="2014-01-01" gender="F" lastname="Popp" firstname="Lotte" license="511994" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:55.85" heatid="3005" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:44.81" heatid="7010" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:00.00" heatid="13001" lane="1" />
                <ENTRY eventid="15" entrytime="00:00:00.00" heatid="15001" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:44.96" heatid="19006" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2135" eventid="3" swimtime="00:00:52.40" lane="2" heatid="3005" points="111" />
                <RESULT resultid="2136" eventid="7" swimtime="00:00:45.21" lane="3" heatid="7010" points="130" />
                <RESULT resultid="2137" eventid="13" swimtime="00:00:50.92" lane="1" heatid="13001" points="109" />
                <RESULT resultid="2138" eventid="15" swimtime="00:02:02.07" lane="1" heatid="15001" points="90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2139" eventid="19" swimtime="00:01:45.33" lane="2" heatid="19006" points="108">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="466" birthdate="2015-01-01" gender="F" lastname="Preißler" firstname="Amy" license="480947" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:59.38" heatid="3003" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:48.04" heatid="7008" lane="3" />
                <ENTRY eventid="15" entrytime="00:00:00.00" heatid="15002" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:48.74" heatid="19005" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2140" eventid="3" swimtime="00:00:53.30" lane="3" heatid="3003" points="106" />
                <RESULT resultid="2141" eventid="7" swimtime="00:00:45.06" lane="3" heatid="7008" points="131" />
                <RESULT resultid="2142" eventid="15" swimtime="00:02:00.57" lane="3" heatid="15002" points="94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2143" eventid="19" swimtime="00:01:46.85" lane="3" heatid="19005" points="104">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="467" birthdate="1992-01-01" gender="F" lastname="Razeto" firstname="Luisa Marie" license="125894" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:25.43" heatid="43000" lane="0" />
                <ENTRY eventid="27" entrytime="00:00:34.07" heatid="27000" lane="0" />
                <ENTRY eventid="41" entrytime="00:00:27.25" heatid="41000" lane="0" />
                <ENTRY eventid="25" entrytime="00:00:28.72" heatid="25000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2144" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
                <RESULT resultid="2145" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="2146" eventid="41" status="WDR" swimtime="00:00:00.00" lane="0" heatid="41000" />
                <RESULT resultid="2147" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="468" birthdate="1986-01-01" gender="M" lastname="Razeto" firstname="Stefano" license="86506" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:21.94" heatid="44017" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:28.42" heatid="28000" lane="0" />
                <ENTRY eventid="42" entrytime="00:00:23.51" heatid="42013" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:24.48" heatid="26010" lane="2" />
                <ENTRY eventid="70" entrytime="00:00:22.36" heatid="70001" lane="2" />
                <ENTRY eventid="66" entrytime="00:00:24.25" heatid="66001" lane="2" />
                <ENTRY eventid="58" entrytime="00:00:25.92" heatid="58001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2148" eventid="44" swimtime="00:00:22.36" lane="2" heatid="44017" points="732" />
                <RESULT resultid="2149" eventid="28" status="WDR" swimtime="00:00:00.00" lane="0" heatid="28000" />
                <RESULT resultid="2150" eventid="42" swimtime="00:00:24.25" lane="2" heatid="42013" points="721" />
                <RESULT resultid="2151" eventid="26" swimtime="00:00:25.92" lane="2" heatid="26010" points="620" />
                <RESULT resultid="2359" eventid="58" swimtime="00:00:24.67" lane="2" heatid="58001" points="719" />
                <RESULT resultid="2343" eventid="66" swimtime="00:00:23.63" lane="2" heatid="66001" points="779" />
                <RESULT resultid="2311" eventid="70" swimtime="00:00:22.28" lane="2" heatid="70001" points="740" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="469" birthdate="2013-01-01" gender="M" lastname="Rebentrost" firstname="Helios" license="461954" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:33.10" heatid="2002" lane="3" />
                <ENTRY eventid="4" entrytime="00:00:42.85" heatid="4015" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:35.95" heatid="8014" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:32.81" heatid="10005" lane="4" />
                <ENTRY eventid="14" entrytime="00:00:37.61" heatid="14007" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:22.00" heatid="20012" lane="4" />
                <ENTRY eventid="22" entrytime="00:03:30.86" heatid="22002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2152" eventid="2" swimtime="00:01:36.00" lane="3" heatid="2002" points="123">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2153" eventid="4" swimtime="00:00:41.73" lane="4" heatid="4015" points="148" />
                <RESULT resultid="2154" eventid="8" swimtime="00:00:34.03" lane="1" heatid="8014" points="207" />
                <RESULT resultid="2155" eventid="10" swimtime="00:01:28.81" lane="4" heatid="10005" points="170">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2156" eventid="14" swimtime="00:00:37.57" lane="1" heatid="14007" points="194" />
                <RESULT resultid="2157" eventid="20" swimtime="00:01:22.07" lane="4" heatid="20012" points="163">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2158" eventid="22" swimtime="00:03:20.13" lane="1" heatid="22002" points="164">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:34.39" />
                    <SPLIT distance="150" swimtime="00:02:33.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="470" birthdate="2015-01-01" gender="M" lastname="Reuße" firstname="Ben" license="484406" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:56.55" heatid="4002" lane="1" />
                <ENTRY eventid="6" entrytime="00:02:02.54" heatid="6002" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:51.43" heatid="8003" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:53.88" heatid="18005" lane="1" />
                <ENTRY eventid="20" entrytime="00:02:06.46" heatid="20001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2159" eventid="4" swimtime="00:00:56.12" lane="1" heatid="4002" points="61" />
                <RESULT resultid="2160" eventid="6" swimtime="00:02:00.38" lane="2" heatid="6002" points="96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2161" eventid="8" swimtime="00:00:49.17" lane="3" heatid="8003" points="68" />
                <RESULT resultid="2162" eventid="18" swimtime="00:00:56.19" lane="1" heatid="18005" points="87" />
                <RESULT resultid="2163" eventid="20" swimtime="00:01:53.19" lane="3" heatid="20001" points="62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="471" birthdate="2007-01-01" gender="M" lastname="Richter" firstname="Kimi" license="384061" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.90" heatid="44000" lane="0" />
                <ENTRY eventid="28" entrytime="00:00:31.92" heatid="28000" lane="0" />
                <ENTRY eventid="48" entrytime="00:01:03.22" heatid="48000" lane="0" />
                <ENTRY eventid="42" entrytime="00:00:28.00" heatid="42000" lane="0" />
                <ENTRY eventid="26" entrytime="00:00:28.10" heatid="26000" lane="0" />
                <ENTRY eventid="32" entrytime="00:00:55.77" heatid="32000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2164" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="2165" eventid="28" status="WDR" swimtime="00:00:00.00" lane="0" heatid="28000" />
                <RESULT resultid="2166" eventid="48" status="WDR" swimtime="00:00:00.00" lane="0" heatid="48000" />
                <RESULT resultid="2167" eventid="42" status="WDR" swimtime="00:00:00.00" lane="0" heatid="42000" />
                <RESULT resultid="2168" eventid="26" status="WDR" swimtime="00:00:00.00" lane="0" heatid="26000" />
                <RESULT resultid="2169" eventid="32" status="WDR" swimtime="00:00:00.00" lane="0" heatid="32000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="472" birthdate="2002-01-01" gender="F" lastname="Richter" firstname="Nele" license="402475" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:28.89" heatid="43014" lane="2" />
                <ENTRY eventid="29" entrytime="00:01:11.85" heatid="29006" lane="4" />
                <ENTRY eventid="51" entrytime="00:02:26.36" heatid="51002" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:30.96" heatid="41012" lane="2" />
                <ENTRY eventid="25" entrytime="00:00:32.66" heatid="25009" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:03.27" heatid="31013" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2170" eventid="43" swimtime="00:00:28.48" lane="2" heatid="43014" points="521" />
                <RESULT resultid="2171" eventid="29" swimtime="00:01:12.31" lane="4" heatid="29006" points="417">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2172" eventid="51" swimtime="00:02:28.23" lane="3" heatid="51002" points="412">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:08.30" />
                    <SPLIT distance="150" swimtime="00:01:48.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2173" eventid="41" swimtime="00:00:31.57" lane="2" heatid="41012" points="460" />
                <RESULT resultid="2174" eventid="25" swimtime="00:00:33.01" lane="2" heatid="25009" points="447" />
                <RESULT resultid="2175" eventid="31" swimtime="00:01:05.95" lane="2" heatid="31013" points="442">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="473" birthdate="2008-01-01" gender="F" lastname="Richter" firstname="Tine" license="429666" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.81" heatid="43013" lane="1" />
                <ENTRY eventid="29" entrytime="00:01:22.03" heatid="29006" lane="1" />
                <ENTRY eventid="47" entrytime="00:01:20.90" heatid="47007" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:33.63" heatid="41011" lane="1" />
                <ENTRY eventid="25" entrytime="00:00:35.81" heatid="25008" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:09.46" heatid="31012" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2176" eventid="43" swimtime="00:00:30.51" lane="1" heatid="43013" points="424" />
                <RESULT resultid="2177" eventid="29" swimtime="00:01:20.71" lane="1" heatid="29006" points="300">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2178" eventid="47" swimtime="00:01:20.89" lane="1" heatid="47007" points="312">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2179" eventid="41" swimtime="00:00:33.64" lane="1" heatid="41011" points="380" />
                <RESULT resultid="2180" eventid="25" swimtime="00:00:36.73" lane="3" heatid="25008" points="324" />
                <RESULT resultid="2181" eventid="31" swimtime="00:01:11.67" lane="4" heatid="31012" points="344">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="474" birthdate="2011-01-01" gender="F" lastname="Rößler" firstname="Lina" license="476556" nation="GER">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:47.46" heatid="27001" lane="1" />
                <ENTRY eventid="47" entrytime="00:01:40.00" heatid="47001" lane="1" />
                <ENTRY eventid="33" entrytime="00:01:39.57" heatid="33001" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:43.57" heatid="41001" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:43.61" heatid="25001" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:49.03" heatid="45001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2182" eventid="27" swimtime="00:00:47.32" lane="1" heatid="27001" points="215" />
                <RESULT resultid="2183" eventid="47" swimtime="00:01:41.12" lane="1" heatid="47001" points="159">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2184" eventid="33" swimtime="00:01:37.20" lane="3" heatid="33001" points="196">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2185" eventid="41" swimtime="00:00:42.05" lane="3" heatid="41001" points="194" />
                <RESULT resultid="2186" eventid="25" swimtime="00:00:45.07" lane="2" heatid="25001" points="175" />
                <RESULT resultid="2187" eventid="45" swimtime="00:01:43.00" lane="1" heatid="45001" points="221">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="475" birthdate="2015-01-01" gender="F" lastname="Sachse" firstname="Luna" license="497634" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:59.16" heatid="3004" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:50.62" heatid="7006" lane="3" />
                <ENTRY eventid="15" entrytime="00:00:00.00" heatid="15001" lane="3" />
                <ENTRY eventid="19" entrytime="00:02:10.39" heatid="19002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2188" eventid="3" swimtime="00:00:53.69" lane="4" heatid="3004" points="104" />
                <RESULT resultid="2189" eventid="7" swimtime="00:00:49.81" lane="3" heatid="7006" points="97" />
                <RESULT resultid="2190" eventid="15" swimtime="00:02:01.74" lane="3" heatid="15001" points="91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2191" eventid="19" swimtime="00:02:07.66" lane="1" heatid="19002" points="60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="478" birthdate="2011-01-01" gender="F" lastname="Schreiter" firstname="Melissa" license="447078" nation="GER">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:36.67" heatid="27000" lane="0" />
                <ENTRY eventid="47" entrytime="00:01:17.50" heatid="47000" lane="0" />
                <ENTRY eventid="37" entrytime="00:02:46.59" heatid="37000" lane="0" />
                <ENTRY eventid="25" entrytime="00:00:34.82" heatid="25000" lane="0" />
                <ENTRY eventid="45" entrytime="00:01:18.35" heatid="45000" lane="0" />
                <ENTRY eventid="53" entrytime="00:02:35.18" heatid="53000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2199" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="2200" eventid="47" status="WDR" swimtime="00:00:00.00" lane="0" heatid="47000" />
                <RESULT resultid="2201" eventid="37" status="WDR" swimtime="00:00:00.00" lane="0" heatid="37000" />
                <RESULT resultid="2202" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
                <RESULT resultid="2203" eventid="45" status="WDR" swimtime="00:00:00.00" lane="0" heatid="45000" />
                <RESULT resultid="2204" eventid="53" status="WDR" swimtime="00:00:00.00" lane="0" heatid="53000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="479" birthdate="2010-01-01" gender="M" lastname="Schrepel" firstname="Alois" license="461950" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:33.83" heatid="44002" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:45.05" heatid="28001" lane="3" />
                <ENTRY eventid="34" entrytime="00:01:38.05" heatid="34001" lane="1" />
                <ENTRY eventid="52" entrytime="00:03:02.36" heatid="52001" lane="2" />
                <ENTRY eventid="46" entrytime="00:01:43.40" heatid="46001" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:23.62" heatid="32001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2205" eventid="44" swimtime="00:00:32.07" lane="1" heatid="44002" points="248" />
                <RESULT resultid="2206" eventid="28" swimtime="00:00:43.58" lane="3" heatid="28001" points="187" />
                <RESULT resultid="2207" eventid="34" status="DSQ" swimtime="00:01:28.56" lane="1" heatid="34001" comment="Der Sportler startete vor dem Startsignal">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2208" eventid="52" swimtime="00:02:59.58" lane="2" heatid="52001" points="169">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:27.09" />
                    <SPLIT distance="150" swimtime="00:02:16.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2209" eventid="46" swimtime="00:01:41.62" lane="4" heatid="46001" points="160">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2210" eventid="32" swimtime="00:01:19.43" lane="1" heatid="32001" points="179">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="480" birthdate="2007-01-01" gender="M" lastname="Schrepel" firstname="Johannes" license="393375" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:28.73" heatid="44000" lane="0" />
                <ENTRY eventid="28" entrytime="00:00:36.46" heatid="28000" lane="0" />
                <ENTRY eventid="42" entrytime="00:00:32.57" heatid="42000" lane="0" />
                <ENTRY eventid="26" entrytime="00:00:34.21" heatid="26000" lane="0" />
                <ENTRY eventid="32" entrytime="00:01:05.69" heatid="32000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2211" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="2212" eventid="28" status="WDR" swimtime="00:00:00.00" lane="0" heatid="28000" />
                <RESULT resultid="2213" eventid="42" status="WDR" swimtime="00:00:00.00" lane="0" heatid="42000" />
                <RESULT resultid="2214" eventid="26" status="WDR" swimtime="00:00:00.00" lane="0" heatid="26000" />
                <RESULT resultid="2215" eventid="32" status="WDR" swimtime="00:00:00.00" lane="0" heatid="32000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="481" birthdate="2014-01-01" gender="M" lastname="Steiner" firstname="Alexander B." license="458124" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:02:01.29" heatid="2001" lane="4" />
                <ENTRY eventid="6" entrytime="00:01:49.58" heatid="6004" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:42.36" heatid="8008" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:51.85" heatid="14002" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:49.23" heatid="18006" lane="2" />
                <ENTRY eventid="38" entrytime="00:04:09.49" heatid="38001" lane="1" />
                <ENTRY eventid="50" entrytime="00:04:36.66" heatid="50001" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:41.67" heatid="20004" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2216" eventid="2" swimtime="00:02:02.68" lane="4" heatid="2001" points="59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2217" eventid="6" swimtime="00:01:47.80" lane="1" heatid="6004" points="134">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2218" eventid="8" swimtime="00:00:41.89" lane="3" heatid="8008" points="111" />
                <RESULT resultid="2219" eventid="14" swimtime="00:00:58.13" lane="2" heatid="14002" points="52" />
                <RESULT resultid="2220" eventid="18" swimtime="00:00:50.03" lane="2" heatid="18006" points="124" />
                <RESULT resultid="2294" eventid="20" swimtime="00:01:44.08" lane="1" heatid="20004" points="79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2221" eventid="38" swimtime="00:04:03.98" lane="1" heatid="38001" points="119">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.04" />
                    <SPLIT distance="100" swimtime="00:01:56.45" />
                    <SPLIT distance="150" swimtime="00:03:02.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2222" eventid="50" swimtime="00:04:40.19" lane="3" heatid="50001" points="55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.51" />
                    <SPLIT distance="100" swimtime="00:02:12.29" />
                    <SPLIT distance="150" swimtime="00:03:29.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="482" birthdate="2013-01-01" gender="F" lastname="Steinert" firstname="Charlotte" license="497631" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:47.31" heatid="3012" lane="4" />
                <ENTRY eventid="5" entrytime="00:01:57.32" heatid="5004" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:41.63" heatid="7014" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:46.20" heatid="15007" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:51.26" heatid="17010" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:32.53" heatid="19012" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2223" eventid="3" status="DSQ" swimtime="00:00:46.11" lane="4" heatid="3012" comment="Die Sportlerin startete vor dem Startsignal" />
                <RESULT resultid="2224" eventid="5" swimtime="00:01:48.76" lane="3" heatid="5004" points="188">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2225" eventid="7" swimtime="00:00:39.65" lane="1" heatid="7014" points="193" />
                <RESULT resultid="2226" eventid="15" swimtime="00:01:43.36" lane="2" heatid="15007" points="149">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2227" eventid="17" swimtime="00:00:51.81" lane="1" heatid="17010" points="164" />
                <RESULT resultid="2228" eventid="19" swimtime="00:01:32.55" lane="1" heatid="19012" points="160">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="483" birthdate="2013-01-01" gender="F" lastname="Stieglitz" firstname="Zoe" license="480944" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:42.46" heatid="3017" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:36.87" heatid="7020" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:35.99" heatid="9008" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:51.48" heatid="13003" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:34.23" heatid="15012" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:49.55" heatid="17011" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:23.46" heatid="19017" lane="1" />
                <ENTRY eventid="51" entrytime="00:03:09.99" heatid="51001" lane="4" />
                <ENTRY eventid="35" entrytime="00:03:17.43" heatid="35001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2229" eventid="3" swimtime="00:00:40.90" lane="1" heatid="3017" points="235" />
                <RESULT resultid="2230" eventid="7" swimtime="00:00:37.03" lane="3" heatid="7020" points="237" />
                <RESULT resultid="2231" eventid="9" swimtime="00:01:30.04" lane="2" heatid="9008" points="247">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2232" eventid="13" swimtime="00:00:43.04" lane="3" heatid="13003" points="181" />
                <RESULT resultid="2233" eventid="15" swimtime="00:01:33.38" lane="1" heatid="15012" points="203">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2234" eventid="17" swimtime="00:00:48.10" lane="1" heatid="17011" points="205" />
                <RESULT resultid="2235" eventid="19" swimtime="00:01:25.52" lane="1" heatid="19017" points="202">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2236" eventid="51" status="DNS" swimtime="00:00:00.00" lane="4" heatid="51001" />
                <RESULT resultid="2237" eventid="35" status="DNS" swimtime="00:00:00.00" lane="3" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="485" birthdate="2009-01-01" gender="M" lastname="Tutzschky" firstname="Lukas" license="461949" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:28.96" heatid="44006" lane="4" />
                <ENTRY eventid="30" entrytime="00:01:13.66" heatid="30001" lane="2" />
                <ENTRY eventid="48" entrytime="00:01:16.47" heatid="48002" lane="3" />
                <ENTRY eventid="52" entrytime="00:02:20.31" heatid="52004" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:32.15" heatid="42004" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:32.87" heatid="26004" lane="2" />
                <ENTRY eventid="32" entrytime="00:01:02.26" heatid="32005" lane="2" />
                <ENTRY eventid="54" entrytime="00:03:27.91" heatid="54001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2242" eventid="44" swimtime="00:00:27.69" lane="4" heatid="44006" points="385" />
                <RESULT resultid="2243" eventid="30" swimtime="00:01:10.58" lane="2" heatid="30001" points="310">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2244" eventid="48" swimtime="00:01:15.95" lane="3" heatid="48002" points="257">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2245" eventid="52" swimtime="00:02:22.90" lane="1" heatid="52004" points="336">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:50.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2246" eventid="42" swimtime="00:00:31.28" lane="4" heatid="42004" points="336" />
                <RESULT resultid="2247" eventid="26" swimtime="00:00:32.43" lane="2" heatid="26004" points="316" />
                <RESULT resultid="2248" eventid="32" swimtime="00:01:03.65" lane="2" heatid="32005" points="349">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2249" eventid="54" swimtime="00:02:44.05" lane="1" heatid="54001" points="298">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:20.07" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="486" birthdate="2015-01-01" gender="M" lastname="Unger" firstname="Bruno" license="471531" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:33.40" heatid="6009" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:34.31" heatid="8022" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:30.98" heatid="10010" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:42.79" heatid="14009" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:42.93" heatid="18012" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:22.32" heatid="20011" lane="2" />
                <ENTRY eventid="38" entrytime="00:03:38.70" heatid="38002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2250" eventid="6" swimtime="00:01:31.49" lane="3" heatid="6009" points="220">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2251" eventid="8" swimtime="00:00:33.79" lane="2" heatid="8022" points="212" />
                <RESULT resultid="2252" eventid="10" swimtime="00:01:30.95" lane="1" heatid="10010" points="159">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2253" eventid="14" swimtime="00:00:41.33" lane="3" heatid="14009" points="145" />
                <RESULT resultid="2254" eventid="18" swimtime="00:00:41.68" lane="3" heatid="18012" points="214" />
                <RESULT resultid="2255" eventid="20" swimtime="00:01:23.29" lane="2" heatid="20011" points="156">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2256" eventid="38" swimtime="00:03:21.13" lane="3" heatid="38002" points="213">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:38.04" />
                    <SPLIT distance="150" swimtime="00:02:31.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="487" birthdate="2017-01-01" gender="F" lastname="Unger" firstname="Sonja" license="508118" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:02:01.05" heatid="5011" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:51.52" heatid="7005" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:52.47" heatid="17016" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2257" eventid="5" swimtime="00:01:55.70" lane="3" heatid="5011" points="156">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2258" eventid="7" swimtime="00:00:53.81" lane="3" heatid="7005" points="77" />
                <RESULT resultid="2259" eventid="17" swimtime="00:00:51.83" lane="2" heatid="17016" points="163" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="490" birthdate="2005-01-01" gender="M" lastname="Weiß" firstname="Johann" license="327133" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:28.32" heatid="44006" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:33.23" heatid="28007" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2266" eventid="44" swimtime="00:00:27.83" lane="2" heatid="44006" points="380" />
                <RESULT resultid="2267" eventid="28" swimtime="00:00:33.92" lane="4" heatid="28007" points="397" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="491" birthdate="2002-01-01" gender="M" lastname="Weiß" firstname="Konrad" license="298099" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:28.21" heatid="44007" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:36.02" heatid="28005" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2268" eventid="44" swimtime="00:00:29.97" lane="4" heatid="44007" points="304" />
                <RESULT resultid="2269" eventid="28" swimtime="00:00:38.25" lane="4" heatid="28005" points="277" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="492" birthdate="1994-01-01" gender="M" lastname="Wewetzer" firstname="Frederik" license="247404" nation="GER">
              <ENTRIES>
                <ENTRY eventid="32" entrytime="00:01:02.59" heatid="32000" lane="0" />
                <ENTRY eventid="44" entrytime="00:00:28.16" heatid="44000" lane="0" />
                <ENTRY eventid="28" entrytime="00:00:34.67" heatid="28000" lane="0" />
                <ENTRY eventid="46" entrytime="00:01:17.36" heatid="46000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2270" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="2271" eventid="28" status="WDR" swimtime="00:00:00.00" lane="0" heatid="28000" />
                <RESULT resultid="2272" eventid="46" status="WDR" swimtime="00:00:00.00" lane="0" heatid="46000" />
                <RESULT resultid="2273" eventid="32" status="WDR" swimtime="00:00:00.00" lane="0" heatid="32000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="497" birthdate="2011-01-01" gender="M" lastname="Britsche" firstname="Jamie Joel" license="0" nation="GER">
              <ENTRIES>
                <ENTRY eventid="26" entrytime="00:00:00.00" heatid="26001" lane="4" />
                <ENTRY eventid="44" entrytime="00:00:00.00" heatid="44001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2295" eventid="44" swimtime="00:00:41.87" lane="4" heatid="44001" points="111" />
                <RESULT resultid="2297" eventid="26" swimtime="00:00:44.35" lane="4" heatid="26001" points="123" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:49.99" lane="3" heatid="40002" />
                <ENTRY eventid="72" entrytime="00:01:59.99" lane="3" heatid="72002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1845" eventid="40" swimtime="00:01:44.79" lane="3" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.23" />
                    <SPLIT distance="100" swimtime="00:00:49.61" />
                    <SPLIT distance="150" swimtime="00:01:16.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="468" number="1" />
                    <RELAYPOSITION athleteid="459" number="2" />
                    <RELAYPOSITION athleteid="485" number="3" />
                    <RELAYPOSITION athleteid="490" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1846" eventid="72" swimtime="00:01:55.34" lane="3" heatid="72002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.13" />
                    <SPLIT distance="100" swimtime="00:00:57.90" />
                    <SPLIT distance="150" swimtime="00:01:28.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="468" number="1" />
                    <RELAYPOSITION athleteid="490" number="2" />
                    <RELAYPOSITION athleteid="425" number="3" />
                    <RELAYPOSITION athleteid="485" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:02:02.39" lane="1" heatid="39002" />
                <ENTRY eventid="71" entrytime="00:02:14.56" lane="3" heatid="71002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1847" eventid="39" swimtime="00:02:02.22" lane="1" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="100" swimtime="00:00:59.22" />
                    <SPLIT distance="150" swimtime="00:01:30.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="472" number="1" />
                    <RELAYPOSITION athleteid="473" number="2" />
                    <RELAYPOSITION athleteid="457" number="3" />
                    <RELAYPOSITION athleteid="434" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1848" eventid="71" swimtime="00:02:16.48" lane="3" heatid="71002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:45.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="472" number="1" />
                    <RELAYPOSITION athleteid="439" number="2" />
                    <RELAYPOSITION athleteid="473" number="3" />
                    <RELAYPOSITION athleteid="457" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:09.99" lane="4" heatid="11003" />
                <ENTRY eventid="23" entrytime="00:02:24.99" lane="2" heatid="23002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1849" eventid="11" swimtime="00:02:10.83" lane="4" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:03.41" />
                    <SPLIT distance="150" swimtime="00:01:37.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="454" number="1" />
                    <RELAYPOSITION athleteid="422" number="2" />
                    <RELAYPOSITION athleteid="469" number="3" />
                    <RELAYPOSITION athleteid="463" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1850" eventid="23" swimtime="00:02:31.15" lane="2" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:01:56.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="454" number="1" />
                    <RELAYPOSITION athleteid="446" number="2" />
                    <RELAYPOSITION athleteid="469" number="3" />
                    <RELAYPOSITION athleteid="463" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:54.99" lane="4" heatid="40002" />
                <ENTRY eventid="72" entrytime="00:02:09.99" lane="4" heatid="72002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1851" eventid="40" swimtime="00:01:58.20" lane="4" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="100" swimtime="00:00:58.05" />
                    <SPLIT distance="150" swimtime="00:01:28.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="425" number="1" />
                    <RELAYPOSITION athleteid="491" number="2" />
                    <RELAYPOSITION athleteid="432" number="3" />
                    <RELAYPOSITION athleteid="447" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1852" eventid="72" swimtime="00:02:12.92" lane="4" heatid="72002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:12.25" />
                    <SPLIT distance="150" swimtime="00:01:42.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="447" number="1" />
                    <RELAYPOSITION athleteid="432" number="2" />
                    <RELAYPOSITION athleteid="459" number="3" />
                    <RELAYPOSITION athleteid="491" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:02:04.99" lane="3" heatid="39001" />
                <ENTRY eventid="71" entrytime="00:02:19.99" lane="2" heatid="71001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1853" eventid="39" swimtime="00:02:15.77" lane="3" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:41.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="439" number="1" />
                    <RELAYPOSITION athleteid="458" number="2" />
                    <RELAYPOSITION athleteid="463" number="3" />
                    <RELAYPOSITION athleteid="452" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1854" eventid="71" swimtime="00:02:31.45" lane="2" heatid="71001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="150" swimtime="00:01:56.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="434" number="1" />
                    <RELAYPOSITION athleteid="449" number="2" />
                    <RELAYPOSITION athleteid="458" number="3" />
                    <RELAYPOSITION athleteid="463" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:19.99" lane="4" heatid="11002" />
                <ENTRY eventid="23" entrytime="00:02:34.99" lane="3" heatid="23002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1855" eventid="11" swimtime="00:02:19.32" lane="4" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:43.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="446" number="1" />
                    <RELAYPOSITION athleteid="430" number="2" />
                    <RELAYPOSITION athleteid="450" number="3" />
                    <RELAYPOSITION athleteid="445" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1856" eventid="23" swimtime="00:02:40.54" lane="3" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:04.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="422" number="1" />
                    <RELAYPOSITION athleteid="450" number="2" />
                    <RELAYPOSITION athleteid="483" number="3" />
                    <RELAYPOSITION athleteid="431" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:02:09.99" lane="3" heatid="40001" />
                <ENTRY eventid="72" entrytime="00:02:29.99" lane="2" heatid="72001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1857" eventid="40" swimtime="00:02:10.57" lane="3" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="150" swimtime="00:01:39.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="479" number="1" />
                    <RELAYPOSITION athleteid="423" number="2" />
                    <RELAYPOSITION athleteid="427" number="3" />
                    <RELAYPOSITION athleteid="454" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1858" eventid="72" swimtime="00:02:31.36" lane="2" heatid="72001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:01:58.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="427" number="1" />
                    <RELAYPOSITION athleteid="486" number="2" />
                    <RELAYPOSITION athleteid="423" number="3" />
                    <RELAYPOSITION athleteid="479" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:02:14.99" lane="1" heatid="39001" />
                <ENTRY eventid="71" entrytime="00:02:34.99" lane="3" heatid="71001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1859" eventid="39" swimtime="00:02:37.93" lane="1" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:01:56.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="449" number="1" />
                    <RELAYPOSITION athleteid="462" number="2" />
                    <RELAYPOSITION athleteid="474" number="3" />
                    <RELAYPOSITION athleteid="460" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1860" eventid="71" swimtime="00:02:48.97" lane="3" heatid="71001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:30.18" />
                    <SPLIT distance="150" swimtime="00:02:09.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="474" number="1" />
                    <RELAYPOSITION athleteid="445" number="2" />
                    <RELAYPOSITION athleteid="452" number="3" />
                    <RELAYPOSITION athleteid="460" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:29.99" lane="2" heatid="11001" />
                <ENTRY eventid="23" entrytime="00:02:44.99" lane="1" heatid="23002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1861" eventid="11" swimtime="00:02:28.80" lane="2" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:12.47" />
                    <SPLIT distance="150" swimtime="00:01:48.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="435" number="1" />
                    <RELAYPOSITION athleteid="483" number="2" />
                    <RELAYPOSITION athleteid="431" number="3" />
                    <RELAYPOSITION athleteid="482" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1862" eventid="23" swimtime="00:02:55.27" lane="1" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="100" swimtime="00:01:29.96" />
                    <SPLIT distance="150" swimtime="00:02:14.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="430" number="1" />
                    <RELAYPOSITION athleteid="435" number="2" />
                    <RELAYPOSITION athleteid="445" number="3" />
                    <RELAYPOSITION athleteid="482" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="72" entrytime="00:02:39.99" lane="3" heatid="72001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1863" eventid="72" status="DNS" swimtime="00:00:00.00" lane="3" heatid="72001" />
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="71" entrytime="00:02:44.99" lane="1" heatid="71001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1864" eventid="71" status="DNS" swimtime="00:00:00.00" lane="1" heatid="71001" />
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:39.99" lane="3" heatid="11001" />
                <ENTRY eventid="23" entrytime="00:02:59.99" lane="2" heatid="23001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1865" eventid="11" swimtime="00:02:48.29" lane="3" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:05.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="481" number="1" />
                    <RELAYPOSITION athleteid="451" number="2" />
                    <RELAYPOSITION athleteid="428" number="3" />
                    <RELAYPOSITION athleteid="437" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1866" eventid="23" swimtime="00:02:58.79" lane="2" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                    <SPLIT distance="100" swimtime="00:01:29.35" />
                    <SPLIT distance="150" swimtime="00:02:20.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="428" number="1" />
                    <RELAYPOSITION athleteid="424" number="2" />
                    <RELAYPOSITION athleteid="481" number="3" />
                    <RELAYPOSITION athleteid="451" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SV 1919 Grimma" nation="GER" region="12" code="5149">
          <ATHLETES>
            <ATHLETE athleteid="71" birthdate="2014-01-01" gender="M" lastname="Adler" firstname="Matteo" license="451964">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:42.75" heatid="2003" lane="1" />
                <ENTRY eventid="4" entrytime="00:00:40.27" heatid="4010" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:33.48" heatid="8017" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:30.69" heatid="10005" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:42.56" heatid="14005" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:17.23" heatid="20013" lane="1" />
                <ENTRY eventid="22" entrytime="00:03:32.67" heatid="22003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="285" eventid="2" swimtime="00:01:39.02" lane="1" heatid="2003" points="112">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="286" eventid="4" swimtime="00:00:38.97" lane="2" heatid="4010" points="182" />
                <RESULT resultid="287" eventid="8" swimtime="00:00:32.87" lane="2" heatid="8017" points="230" />
                <RESULT resultid="288" eventid="10" swimtime="00:01:28.51" lane="2" heatid="10005" points="172">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="289" eventid="14" swimtime="00:00:44.24" lane="1" heatid="14005" points="118" />
                <RESULT resultid="290" eventid="20" swimtime="00:01:17.37" lane="1" heatid="20013" points="194">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="291" eventid="22" swimtime="00:03:14.48" lane="1" heatid="22003" points="179">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:34.18" />
                    <SPLIT distance="150" swimtime="00:02:33.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="72" birthdate="2015-01-01" gender="M" lastname="Anders" firstname="Erwin Max" license="482472">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:47.02" heatid="4013" lane="1" />
                <ENTRY eventid="6" entrytime="00:01:45.99" heatid="6005" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:36.92" heatid="8012" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:43.97" heatid="16008" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:48.56" heatid="18012" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:24.86" heatid="20010" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="292" eventid="4" swimtime="00:00:45.61" lane="1" heatid="4013" points="113" />
                <RESULT resultid="293" eventid="6" swimtime="00:01:46.53" lane="4" heatid="6005" points="139">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="294" eventid="8" status="DNS" swimtime="00:00:00.00" lane="3" heatid="8012" />
                <RESULT resultid="295" eventid="16" swimtime="00:01:39.22" lane="1" heatid="16008" points="115">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="296" eventid="18" swimtime="00:00:50.34" lane="4" heatid="18012" points="121" />
                <RESULT resultid="297" eventid="20" swimtime="00:01:21.92" lane="3" heatid="20010" points="163">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="73" birthdate="2015-01-01" gender="F" lastname="Dozsa-Nemeth" firstname="Odett" license="463478">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:38.73" heatid="3021" lane="2" />
                <ENTRY eventid="5" entrytime="00:01:41.46" heatid="5013" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:35.46" heatid="7028" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:25.78" heatid="15017" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:46.57" heatid="17018" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:23.58" heatid="19017" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="298" eventid="3" swimtime="00:00:37.70" lane="2" heatid="3021" points="300" />
                <RESULT resultid="299" eventid="5" swimtime="00:01:41.39" lane="1" heatid="5013" points="232">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="300" eventid="7" swimtime="00:00:35.81" lane="4" heatid="7028" points="262" />
                <RESULT resultid="301" eventid="15" swimtime="00:01:22.55" lane="3" heatid="15017" points="293">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="302" eventid="17" swimtime="00:00:47.03" lane="1" heatid="17018" points="219" />
                <RESULT resultid="303" eventid="19" swimtime="00:01:24.92" lane="4" heatid="19017" points="207">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="74" birthdate="2010-01-01" gender="M" lastname="Duckstein" firstname="Alex" license="412300">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:28.23" heatid="44000" lane="0" />
                <ENTRY eventid="28" entrytime="00:00:37.05" heatid="28000" lane="0" />
                <ENTRY eventid="48" entrytime="00:01:15.79" heatid="48000" lane="0" />
                <ENTRY eventid="34" entrytime="00:01:12.71" heatid="34000" lane="0" />
                <ENTRY eventid="42" entrytime="00:00:31.12" heatid="42000" lane="0" />
                <ENTRY eventid="26" entrytime="00:00:34.42" heatid="26000" lane="0" />
                <ENTRY eventid="46" entrytime="00:01:27.43" heatid="46000" lane="0" />
                <ENTRY eventid="32" entrytime="00:01:04.37" heatid="32000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="304" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="305" eventid="28" status="WDR" swimtime="00:00:00.00" lane="0" heatid="28000" />
                <RESULT resultid="306" eventid="48" status="WDR" swimtime="00:00:00.00" lane="0" heatid="48000" />
                <RESULT resultid="307" eventid="34" status="WDR" swimtime="00:00:00.00" lane="0" heatid="34000" />
                <RESULT resultid="308" eventid="42" status="WDR" swimtime="00:00:00.00" lane="0" heatid="42000" />
                <RESULT resultid="309" eventid="26" status="WDR" swimtime="00:00:00.00" lane="0" heatid="26000" />
                <RESULT resultid="310" eventid="46" status="WDR" swimtime="00:00:00.00" lane="0" heatid="46000" />
                <RESULT resultid="311" eventid="32" status="WDR" swimtime="00:00:00.00" lane="0" heatid="32000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="75" birthdate="2017-01-01" gender="F" lastname="Gerke" firstname="Lilly" license="501087">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:01:03.98" heatid="3001" lane="2" />
                <ENTRY eventid="5" entrytime="00:02:19.85" heatid="5002" lane="3" />
                <ENTRY eventid="7" entrytime="00:01:01.81" heatid="7001" lane="3" />
                <ENTRY eventid="17" entrytime="00:01:06.50" heatid="17003" lane="2" />
                <ENTRY eventid="19" entrytime="00:02:03.35" heatid="19003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="312" eventid="3" swimtime="00:00:56.62" lane="2" heatid="3001" points="88" />
                <RESULT resultid="313" eventid="5" swimtime="00:02:14.44" lane="3" heatid="5002" points="99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="314" eventid="7" swimtime="00:00:51.09" lane="3" heatid="7001" points="90" />
                <RESULT resultid="315" eventid="17" swimtime="00:01:03.43" lane="2" heatid="17003" points="89" />
                <RESULT resultid="316" eventid="19" swimtime="00:01:56.94" lane="4" heatid="19003" points="79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="76" birthdate="2015-01-01" gender="F" lastname="Golze" firstname="Clara" license="463479">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.20" heatid="3015" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:39.93" heatid="7016" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:45.20" heatid="9005" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:48.27" heatid="13005" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:40.01" heatid="15009" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="317" eventid="3" swimtime="00:00:45.30" lane="1" heatid="3015" points="173" />
                <RESULT resultid="318" eventid="7" swimtime="00:00:40.63" lane="2" heatid="7016" points="179" />
                <RESULT resultid="319" eventid="9" swimtime="00:01:44.79" lane="4" heatid="9005" points="156">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="320" eventid="13" swimtime="00:00:47.77" lane="1" heatid="13005" points="132" />
                <RESULT resultid="321" eventid="15" swimtime="00:01:41.06" lane="3" heatid="15009" points="160">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="77" birthdate="2016-01-01" gender="M" lastname="Haferkorn" firstname="Arne" license="482477">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:45.91" heatid="4012" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:38.22" heatid="8021" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:37.09" heatid="10009" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:47.71" heatid="14008" lane="1" />
                <ENTRY eventid="16" entrytime="00:01:40.95" heatid="16007" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:26.72" heatid="20018" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="322" eventid="4" swimtime="00:00:43.46" lane="1" heatid="4012" points="131" />
                <RESULT resultid="323" eventid="8" swimtime="00:00:37.62" lane="3" heatid="8021" points="153" />
                <RESULT resultid="324" eventid="10" swimtime="00:01:33.91" lane="1" heatid="10009" points="144">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="325" eventid="14" swimtime="00:00:45.28" lane="1" heatid="14008" points="110" />
                <RESULT resultid="326" eventid="16" swimtime="00:01:39.63" lane="1" heatid="16007" points="114">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="327" eventid="20" swimtime="00:01:23.39" lane="3" heatid="20018" points="155">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="78" birthdate="2011-01-01" gender="F" lastname="Harbich" firstname="Svea" license="422683">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.52" heatid="43011" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:41.25" heatid="27007" lane="1" />
                <ENTRY eventid="47" entrytime="00:01:22.36" heatid="47005" lane="3" />
                <ENTRY eventid="25" entrytime="00:00:36.66" heatid="25006" lane="1" />
                <ENTRY eventid="45" entrytime="00:01:29.67" heatid="45005" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:07.94" heatid="31010" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="328" eventid="43" swimtime="00:00:29.93" lane="3" heatid="43011" points="449" />
                <RESULT resultid="329" eventid="27" swimtime="00:00:40.55" lane="1" heatid="27007" points="342" />
                <RESULT resultid="330" eventid="47" swimtime="00:01:19.25" lane="3" heatid="47005" points="332">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="331" eventid="25" swimtime="00:00:36.13" lane="1" heatid="25006" points="341" />
                <RESULT resultid="332" eventid="45" swimtime="00:01:31.00" lane="1" heatid="45005" points="321">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="333" eventid="31" swimtime="00:01:07.40" lane="2" heatid="31010" points="414">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="79" birthdate="2010-01-01" gender="F" lastname="Hartwig" firstname="Annika" license="471349">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:38.39" heatid="27005" lane="1" />
                <ENTRY eventid="29" entrytime="00:01:24.10" heatid="29002" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:22.30" heatid="33004" lane="3" />
                <ENTRY eventid="37" entrytime="00:03:05.67" heatid="37002" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:35.61" heatid="41005" lane="4" />
                <ENTRY eventid="45" entrytime="00:01:23.40" heatid="45006" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:10.30" heatid="31006" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="334" eventid="27" swimtime="00:00:38.53" lane="1" heatid="27005" points="399" />
                <RESULT resultid="335" eventid="29" swimtime="00:01:24.69" lane="3" heatid="29002" points="259">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="336" eventid="33" swimtime="00:01:19.95" lane="3" heatid="33004" points="353">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="337" eventid="37" swimtime="00:03:03.76" lane="4" heatid="37002" points="392">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:01:27.25" />
                    <SPLIT distance="150" swimtime="00:02:15.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="338" eventid="41" swimtime="00:00:35.72" lane="4" heatid="41005" points="317" />
                <RESULT resultid="339" eventid="45" swimtime="00:01:25.52" lane="1" heatid="45006" points="387">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="340" eventid="31" swimtime="00:01:11.16" lane="1" heatid="31006" points="352">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="80" birthdate="2015-01-01" gender="F" lastname="Heinitz" firstname="Linn" license="467472">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:39.23" heatid="5013" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:35.03" heatid="7028" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:32.83" heatid="9011" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:41.18" heatid="13014" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:45.76" heatid="17018" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:20.52" heatid="19023" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="341" eventid="5" swimtime="00:01:37.19" lane="3" heatid="5013" points="264">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="342" eventid="7" swimtime="00:00:34.25" lane="1" heatid="7028" points="300" />
                <RESULT resultid="343" eventid="9" swimtime="00:01:30.64" lane="4" heatid="9011" points="242">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="344" eventid="13" swimtime="00:00:39.74" lane="3" heatid="13014" points="230" />
                <RESULT resultid="345" eventid="17" swimtime="00:00:43.62" lane="3" heatid="17018" points="275" />
                <RESULT resultid="346" eventid="19" swimtime="00:01:18.68" lane="4" heatid="19023" points="260">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="81" birthdate="2014-01-01" gender="F" lastname="Huerta-Stiehl" firstname="Nelly Johanna" license="451404">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:34.46" heatid="5010" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:36.52" heatid="7021" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:37.78" heatid="9007" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:44.08" heatid="17019" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:23.26" heatid="19017" lane="3" />
                <ENTRY eventid="21" entrytime="00:03:24.74" heatid="21001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="347" eventid="5" swimtime="00:01:33.59" lane="2" heatid="5010" points="295">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="348" eventid="7" swimtime="00:00:35.27" lane="3" heatid="7021" points="274" />
                <RESULT resultid="349" eventid="9" swimtime="00:01:32.14" lane="1" heatid="9007" points="230">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="350" eventid="17" swimtime="00:00:43.02" lane="4" heatid="17019" points="286" />
                <RESULT resultid="351" eventid="19" swimtime="00:01:19.47" lane="3" heatid="19017" points="252">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="352" eventid="21" status="DSQ" swimtime="00:03:19.14" lane="3" heatid="21001" comment="Die Sportlerin hat bei der dritten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                    <SPLIT distance="100" swimtime="00:01:36.77" />
                    <SPLIT distance="150" swimtime="00:02:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="82" birthdate="2016-01-01" gender="F" lastname="Kobsik" firstname="Chiara" license="482474">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:43.71" heatid="3020" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:37.78" heatid="7027" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:40.09" heatid="9015" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:50.50" heatid="13004" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:37.38" heatid="15016" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:25.57" heatid="19022" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="353" eventid="3" swimtime="00:00:42.39" lane="2" heatid="3020" points="211" />
                <RESULT resultid="354" eventid="7" swimtime="00:00:36.15" lane="4" heatid="7027" points="255" />
                <RESULT resultid="355" eventid="9" swimtime="00:01:40.83" lane="3" heatid="9015" points="176">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="356" eventid="13" swimtime="00:00:49.59" lane="3" heatid="13004" points="118" />
                <RESULT resultid="357" eventid="15" swimtime="00:01:34.18" lane="2" heatid="15016" points="197">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="358" eventid="19" swimtime="00:01:25.07" lane="1" heatid="19022" points="206">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="83" birthdate="2012-01-01" gender="F" lastname="Kobsik" firstname="Zoe" license="449834">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:29.73" heatid="43010" lane="2" />
                <ENTRY eventid="29" entrytime="00:01:16.37" heatid="29003" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:18.73" heatid="33006" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:31.33" heatid="41008" lane="2" />
                <ENTRY eventid="25" entrytime="00:00:35.31" heatid="25005" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:05.13" heatid="31009" lane="2" />
                <ENTRY eventid="53" entrytime="00:02:51.22" heatid="53002" lane="3" />
                <ENTRY eventid="55" entrytime="00:00:34.61" heatid="55001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="359" eventid="43" swimtime="00:00:30.02" lane="2" heatid="43010" points="445" />
                <RESULT resultid="360" eventid="29" swimtime="00:01:18.64" lane="2" heatid="29003" points="324">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="361" eventid="33" swimtime="00:01:17.32" lane="1" heatid="33006" points="390">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="362" eventid="41" swimtime="00:00:31.91" lane="2" heatid="41008" points="445" />
                <RESULT resultid="363" eventid="25" swimtime="00:00:34.61" lane="3" heatid="25005" points="388" />
                <RESULT resultid="364" eventid="31" swimtime="00:01:07.85" lane="2" heatid="31009" points="406">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="365" eventid="53" swimtime="00:02:49.53" lane="3" heatid="53002" points="371">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:02:09.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2349" eventid="55" swimtime="00:00:33.56" lane="1" heatid="55001" points="425" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="84" birthdate="2016-01-01" gender="M" lastname="Kühne" firstname="Leon Maurice" license="482481">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:46.78" heatid="4012" lane="4" />
                <ENTRY eventid="6" entrytime="00:02:01.44" heatid="6008" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:41.29" heatid="8009" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:53.15" heatid="14008" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:56.78" heatid="18004" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:33.33" heatid="20018" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="366" eventid="4" swimtime="00:00:47.40" lane="4" heatid="4012" points="101" />
                <RESULT resultid="367" eventid="6" swimtime="00:02:05.00" lane="1" heatid="6008" points="86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="368" eventid="8" swimtime="00:00:43.16" lane="3" heatid="8009" points="101" />
                <RESULT resultid="369" eventid="14" swimtime="00:00:52.95" lane="4" heatid="14008" points="69" />
                <RESULT resultid="370" eventid="18" swimtime="00:00:58.55" lane="4" heatid="18004" points="77" />
                <RESULT resultid="371" eventid="20" swimtime="00:01:33.93" lane="1" heatid="20018" points="108">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="85" birthdate="2017-01-01" gender="M" lastname="Lipinski" firstname="Pepe" license="501094">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:01:00.37" heatid="4001" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:55.23" heatid="8002" lane="1" />
                <ENTRY eventid="10" entrytime="00:00:00.00" heatid="10008" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:56.79" heatid="16006" lane="3" />
                <ENTRY eventid="18" entrytime="00:01:02.66" heatid="18010" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="372" eventid="4" swimtime="00:00:56.52" lane="3" heatid="4001" points="59" />
                <RESULT resultid="373" eventid="8" swimtime="00:00:49.70" lane="1" heatid="8002" points="66" />
                <RESULT resultid="374" eventid="10" swimtime="00:01:59.04" lane="3" heatid="10008" points="70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="375" eventid="16" swimtime="00:02:04.79" lane="3" heatid="16006" points="58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="376" eventid="18" swimtime="00:01:00.75" lane="2" heatid="18010" points="69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="86" birthdate="2009-01-01" gender="F" lastname="Maneck" firstname="Amilia" license="398061">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:28.51" heatid="43009" lane="2" />
                <ENTRY eventid="29" entrytime="00:01:12.78" heatid="29005" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:09.28" heatid="47006" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:13.68" heatid="33005" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:30.76" heatid="41010" lane="4" />
                <ENTRY eventid="25" entrytime="00:00:31.59" heatid="25007" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:02.62" heatid="31011" lane="3" />
                <ENTRY eventid="53" entrytime="00:02:45.72" heatid="53002" lane="2" />
                <ENTRY eventid="67" entrytime="00:00:28.37" heatid="67001" lane="2" />
                <ENTRY eventid="63" entrytime="00:00:31.23" heatid="63001" lane="2" />
                <ENTRY eventid="56" entrytime="00:00:32.19" heatid="56001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="377" eventid="43" swimtime="00:00:28.37" lane="2" heatid="43009" points="528" />
                <RESULT resultid="378" eventid="29" swimtime="00:01:12.64" lane="3" heatid="29005" points="411">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="379" eventid="47" swimtime="00:01:10.99" lane="3" heatid="47006" points="462">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="380" eventid="33" swimtime="00:01:13.84" lane="3" heatid="33005" points="448">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="381" eventid="41" swimtime="00:00:31.23" lane="4" heatid="41010" points="475" />
                <RESULT resultid="382" eventid="25" swimtime="00:00:32.19" lane="4" heatid="25007" points="482" />
                <RESULT resultid="383" eventid="31" swimtime="00:01:02.70" lane="3" heatid="31011" points="514">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="384" eventid="53" swimtime="00:02:45.39" lane="2" heatid="53002" points="399">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:02:07.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2354" eventid="56" swimtime="00:00:31.98" lane="4" heatid="56001" points="492" />
                <RESULT resultid="2331" eventid="63" swimtime="00:00:30.84" lane="2" heatid="63001" points="494" />
                <RESULT resultid="2299" eventid="67" swimtime="00:00:28.05" lane="2" heatid="67001" points="546" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="87" birthdate="2007-01-01" gender="M" lastname="Maneck" firstname="Samuel" license="405759">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.37" heatid="44016" lane="3" />
                <ENTRY eventid="30" entrytime="00:01:01.73" heatid="30005" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:03.47" heatid="34008" lane="2" />
                <ENTRY eventid="52" entrytime="00:02:03.24" heatid="52005" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:26.90" heatid="42012" lane="1" />
                <ENTRY eventid="26" entrytime="00:00:29.03" heatid="26006" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:09.59" heatid="46006" lane="3" />
                <ENTRY eventid="32" entrytime="00:00:53.74" heatid="32012" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="385" eventid="44" swimtime="00:00:24.23" lane="3" heatid="44016" points="575" />
                <RESULT resultid="386" eventid="30" swimtime="00:01:01.48" lane="1" heatid="30005" points="469">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="387" eventid="34" swimtime="00:01:08.58" lane="2" heatid="34008" points="371">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="388" eventid="52" swimtime="00:02:02.88" lane="2" heatid="52005" points="528">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="100" swimtime="00:00:57.38" />
                    <SPLIT distance="150" swimtime="00:01:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="389" eventid="42" swimtime="00:00:27.32" lane="1" heatid="42012" points="504" />
                <RESULT resultid="390" eventid="26" swimtime="00:00:29.52" lane="4" heatid="26006" points="420" />
                <RESULT resultid="391" eventid="46" swimtime="00:01:10.74" lane="3" heatid="46006" points="477">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="392" eventid="32" swimtime="00:00:54.95" lane="3" heatid="32012" points="543">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="88" birthdate="2017-01-01" gender="F" lastname="Munari" firstname="Mina" license="501084">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:59.31" heatid="3003" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:54.97" heatid="7004" lane="4" />
                <ENTRY eventid="15" entrytime="00:02:07.51" heatid="15004" lane="4" />
                <ENTRY eventid="17" entrytime="00:01:09.79" heatid="17003" lane="1" />
                <ENTRY eventid="19" entrytime="00:02:00.92" heatid="19003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="393" eventid="3" swimtime="00:00:57.80" lane="2" heatid="3003" points="83" />
                <RESULT resultid="394" eventid="7" swimtime="00:00:54.33" lane="4" heatid="7004" points="75" />
                <RESULT resultid="395" eventid="15" swimtime="00:02:14.45" lane="4" heatid="15004" points="68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="396" eventid="17" swimtime="00:01:10.51" lane="1" heatid="17003" points="65" />
                <RESULT resultid="397" eventid="19" swimtime="00:02:02.73" lane="3" heatid="19003" points="68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="89" birthdate="2015-01-01" gender="F" lastname="Otto" firstname="Pia" license="463476">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:42.75" heatid="3017" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:36.92" heatid="7020" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:35.75" heatid="9009" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:44.02" heatid="13008" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:35.64" heatid="15011" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:21.42" heatid="19019" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="398" eventid="3" status="DNS" swimtime="00:00:00.00" lane="4" heatid="3017" />
                <RESULT resultid="399" eventid="7" status="DNS" swimtime="00:00:00.00" lane="4" heatid="7020" />
                <RESULT resultid="400" eventid="9" status="DNS" swimtime="00:00:00.00" lane="4" heatid="9009" />
                <RESULT resultid="401" eventid="13" status="DNS" swimtime="00:00:00.00" lane="1" heatid="13008" />
                <RESULT resultid="402" eventid="15" status="DNS" swimtime="00:00:00.00" lane="3" heatid="15011" />
                <RESULT resultid="403" eventid="19" status="DNS" swimtime="00:00:00.00" lane="1" heatid="19019" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="90" birthdate="2014-01-01" gender="M" lastname="Polzin" firstname="Franz" license="451411">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:45.12" heatid="6010" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:34.67" heatid="8016" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:32.04" heatid="10005" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:40.83" heatid="14005" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:28.57" heatid="16005" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:46.99" heatid="18013" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:21.17" heatid="20012" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="404" eventid="6" swimtime="00:01:45.65" lane="4" heatid="6010" points="143">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="405" eventid="8" swimtime="00:00:36.29" lane="4" heatid="8016" points="171" />
                <RESULT resultid="406" eventid="10" swimtime="00:01:29.61" lane="1" heatid="10005" points="166">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="407" eventid="14" swimtime="00:00:42.18" lane="2" heatid="14005" points="137" />
                <RESULT resultid="408" eventid="16" swimtime="00:01:26.69" lane="3" heatid="16005" points="173">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="409" eventid="18" swimtime="00:00:49.49" lane="1" heatid="18013" points="128" />
                <RESULT resultid="410" eventid="20" swimtime="00:01:22.11" lane="1" heatid="20012" points="162">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="91" birthdate="2009-01-01" gender="F" lastname="Rasmussen" firstname="Helen" license="398058">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.45" heatid="43007" lane="3" />
                <ENTRY eventid="29" entrytime="00:01:22.36" heatid="29002" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:21.28" heatid="33004" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:34.40" heatid="41005" lane="1" />
                <ENTRY eventid="25" entrytime="00:00:35.68" heatid="25003" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:08.55" heatid="31007" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="411" eventid="43" swimtime="00:00:30.19" lane="3" heatid="43007" points="438" />
                <RESULT resultid="412" eventid="29" swimtime="00:01:21.18" lane="2" heatid="29002" points="295">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="413" eventid="33" swimtime="00:01:20.82" lane="2" heatid="33004" points="341">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="414" eventid="41" swimtime="00:00:33.50" lane="1" heatid="41005" points="385" />
                <RESULT resultid="415" eventid="25" swimtime="00:00:37.88" lane="3" heatid="25003" points="296" />
                <RESULT resultid="416" eventid="31" swimtime="00:01:09.64" lane="2" heatid="31007" points="375">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="92" birthdate="2015-01-01" gender="M" lastname="Schewelew" firstname="Egor" license="463483">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:45.07" heatid="4013" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:35.96" heatid="8014" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:35.40" heatid="10010" lane="4" />
                <ENTRY eventid="14" entrytime="00:00:47.72" heatid="14009" lane="4" />
                <ENTRY eventid="16" entrytime="00:01:35.86" heatid="16008" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:21.32" heatid="20019" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="417" eventid="4" swimtime="00:00:43.71" lane="2" heatid="4013" points="129" />
                <RESULT resultid="418" eventid="8" swimtime="00:00:36.60" lane="4" heatid="8014" points="167" />
                <RESULT resultid="419" eventid="10" swimtime="00:01:37.23" lane="4" heatid="10010" points="130">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="420" eventid="14" swimtime="00:00:46.35" lane="4" heatid="14009" points="103" />
                <RESULT resultid="421" eventid="16" swimtime="00:01:36.80" lane="2" heatid="16008" points="124">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="422" eventid="20" swimtime="00:01:23.70" lane="4" heatid="20019" points="153">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="93" birthdate="2008-01-01" gender="M" lastname="Schmutzer" firstname="Domenik" license="398057">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:25.18" heatid="44012" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:30.51" heatid="28010" lane="2" />
                <ENTRY eventid="48" entrytime="00:01:05.21" heatid="48005" lane="1" />
                <ENTRY eventid="38" entrytime="00:02:36.83" heatid="38005" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:28.62" heatid="42012" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:29.53" heatid="26005" lane="2" />
                <ENTRY eventid="46" entrytime="00:01:08.18" heatid="46006" lane="2" />
                <ENTRY eventid="32" entrytime="00:00:55.73" heatid="32009" lane="2" />
                <ENTRY eventid="62" entrytime="00:00:30.37" heatid="62001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="423" eventid="44" swimtime="00:00:25.20" lane="2" heatid="44012" points="511" />
                <RESULT resultid="424" eventid="28" swimtime="00:00:30.37" lane="2" heatid="28010" points="554" />
                <RESULT resultid="425" eventid="48" swimtime="00:01:05.49" lane="1" heatid="48005" points="401">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="426" eventid="38" swimtime="00:02:34.35" lane="2" heatid="38005" points="471">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="150" swimtime="00:01:53.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="427" eventid="42" swimtime="00:00:28.89" lane="4" heatid="42012" points="426" />
                <RESULT resultid="428" eventid="26" swimtime="00:00:29.99" lane="2" heatid="26005" points="400" />
                <RESULT resultid="429" eventid="46" swimtime="00:01:09.45" lane="2" heatid="46006" points="504">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="430" eventid="32" swimtime="00:00:56.42" lane="2" heatid="32009" points="501">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2329" eventid="62" swimtime="00:00:30.31" lane="1" heatid="62001" points="557" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="94" birthdate="2014-01-01" gender="F" lastname="Seemann" firstname="Emma" license="451406">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:45.34" heatid="1001" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:34.58" heatid="7025" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:31.92" heatid="9011" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:43.14" heatid="13009" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:44.38" heatid="17015" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:21.64" heatid="19019" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="431" eventid="1" status="DSQ" swimtime="00:01:38.51" lane="2" heatid="1001" comment="Beim Anschlag an der Wende hat die Sportlerin nicht mit beiden Händen gleichzeitig angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="432" eventid="7" swimtime="00:00:35.04" lane="1" heatid="7025" points="280" />
                <RESULT resultid="433" eventid="9" swimtime="00:01:30.93" lane="1" heatid="9011" points="240">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="434" eventid="13" swimtime="00:00:41.83" lane="3" heatid="13009" points="197" />
                <RESULT resultid="435" eventid="17" swimtime="00:00:43.88" lane="3" heatid="17015" points="270" />
                <RESULT resultid="436" eventid="19" swimtime="00:01:20.80" lane="4" heatid="19019" points="240">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="95" birthdate="2013-01-01" gender="M" lastname="Thiele" firstname="Henrik" license="451456">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:21.50" heatid="2005" lane="3" />
                <ENTRY eventid="6" entrytime="00:01:22.67" heatid="6011" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:29.17" heatid="8024" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:15.85" heatid="10012" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:32.44" heatid="14011" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:35.62" heatid="18014" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:06.17" heatid="20021" lane="2" />
                <ENTRY eventid="22" entrytime="00:02:46.46" heatid="22005" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="437" eventid="2" swimtime="00:01:15.57" lane="3" heatid="2005" points="252">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="438" eventid="6" swimtime="00:01:24.60" lane="2" heatid="6011" points="278">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="439" eventid="8" swimtime="00:00:29.15" lane="2" heatid="8024" points="330" />
                <RESULT resultid="440" eventid="10" swimtime="00:01:16.73" lane="2" heatid="10012" points="264">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="441" eventid="14" swimtime="00:00:32.52" lane="2" heatid="14011" points="299" />
                <RESULT resultid="442" eventid="18" swimtime="00:00:37.48" lane="2" heatid="18014" points="294" />
                <RESULT resultid="443" eventid="20" swimtime="00:01:06.87" lane="2" heatid="20021" points="301">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="444" eventid="22" swimtime="00:02:46.82" lane="3" heatid="22005" points="283">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="150" swimtime="00:02:10.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="96" birthdate="2008-01-01" gender="M" lastname="Tloczkowski" firstname="Karl-Moritz" license="381054">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.81" heatid="44016" lane="1" />
                <ENTRY eventid="30" entrytime="00:00:59.18" heatid="30005" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:26.47" heatid="42012" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:28.31" heatid="26009" lane="3" />
                <ENTRY eventid="32" entrytime="00:00:54.21" heatid="32012" lane="1" />
                <ENTRY eventid="54" entrytime="00:02:22.00" heatid="54004" lane="4" />
                <ENTRY eventid="69" entrytime="00:00:24.90" heatid="69001" lane="3" />
                <ENTRY eventid="65" entrytime="00:00:26.54" heatid="65001" lane="2" />
                <ENTRY eventid="57" entrytime="00:00:28.46" heatid="57001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="445" eventid="44" swimtime="00:00:24.90" lane="1" heatid="44016" points="530" />
                <RESULT resultid="446" eventid="30" swimtime="00:00:59.30" lane="3" heatid="30005" points="523">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="447" eventid="42" swimtime="00:00:26.54" lane="3" heatid="42012" points="550" />
                <RESULT resultid="448" eventid="26" swimtime="00:00:28.46" lane="3" heatid="26009" points="468" />
                <RESULT resultid="449" eventid="32" swimtime="00:00:55.08" lane="1" heatid="32012" points="539">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="450" eventid="54" swimtime="00:02:22.48" lane="4" heatid="54004" points="455">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:01:06.12" />
                    <SPLIT distance="150" swimtime="00:01:48.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2357" eventid="57" swimtime="00:00:28.38" lane="1" heatid="57001" points="472" />
                <RESULT resultid="2339" eventid="65" swimtime="00:00:26.04" lane="2" heatid="65001" points="582" />
                <RESULT resultid="2308" eventid="69" swimtime="00:00:24.85" lane="3" heatid="69001" points="533" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="97" birthdate="2017-01-01" gender="F" lastname="Vogt" firstname="Alexandra" license="501085">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:52.05" heatid="3009" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:50.37" heatid="7007" lane="4" />
                <ENTRY eventid="9" entrytime="00:02:08.50" heatid="9002" lane="1" />
                <ENTRY eventid="13" entrytime="00:01:01.00" heatid="13002" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:56.68" heatid="15015" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:48.82" heatid="19005" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="451" eventid="3" swimtime="00:00:50.37" lane="4" heatid="3009" points="125" />
                <RESULT resultid="452" eventid="7" swimtime="00:00:47.71" lane="4" heatid="7007" points="111" />
                <RESULT resultid="453" eventid="9" swimtime="00:01:58.63" lane="1" heatid="9002" points="108">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="454" eventid="13" swimtime="00:01:04.95" lane="4" heatid="13002" points="52" />
                <RESULT resultid="455" eventid="15" swimtime="00:01:54.25" lane="4" heatid="15015" points="110">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="456" eventid="19" swimtime="00:01:50.53" lane="1" heatid="19005" points="93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="98" birthdate="2013-01-01" gender="F" lastname="Voigt" firstname="Sophia" license="444104">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:35.33" heatid="3023" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:31.10" heatid="7030" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:23.12" heatid="9018" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:38.16" heatid="13016" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:17.85" heatid="15019" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:08.83" heatid="19025" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="457" eventid="3" swimtime="00:00:34.73" lane="2" heatid="3023" points="384" />
                <RESULT resultid="458" eventid="7" swimtime="00:00:30.81" lane="2" heatid="7030" points="412" />
                <RESULT resultid="459" eventid="9" swimtime="00:01:23.68" lane="1" heatid="9018" points="307">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="460" eventid="13" swimtime="00:00:40.24" lane="4" heatid="13016" points="222" />
                <RESULT resultid="461" eventid="15" swimtime="00:01:18.74" lane="2" heatid="15019" points="338">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="462" eventid="19" swimtime="00:01:08.69" lane="2" heatid="19025" points="391">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="99" birthdate="2005-01-01" gender="M" lastname="von Thun" firstname="Karl" license="329642">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.25" heatid="44013" lane="2" />
                <ENTRY eventid="30" entrytime="00:00:55.29" heatid="30006" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:25.64" heatid="42013" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:26.71" heatid="26010" lane="1" />
                <ENTRY eventid="32" entrytime="00:00:52.06" heatid="32013" lane="3" />
                <ENTRY eventid="70" entrytime="00:00:23.83" heatid="70001" lane="3" />
                <ENTRY eventid="66" entrytime="00:00:25.59" heatid="66001" lane="4" />
                <ENTRY eventid="58" entrytime="00:00:26.64" heatid="58001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="463" eventid="44" swimtime="00:00:23.83" lane="2" heatid="44013" points="605" />
                <RESULT resultid="464" eventid="30" swimtime="00:00:55.12" lane="2" heatid="30006" points="651">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="465" eventid="42" swimtime="00:00:25.59" lane="4" heatid="42013" points="613" />
                <RESULT resultid="466" eventid="26" swimtime="00:00:26.64" lane="1" heatid="26010" points="571" />
                <RESULT resultid="467" eventid="32" swimtime="00:00:51.82" lane="3" heatid="32013" points="647">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2361" eventid="58" swimtime="00:00:26.42" lane="1" heatid="58001" points="586" />
                <RESULT resultid="2346" eventid="66" swimtime="00:00:25.46" lane="4" heatid="66001" points="623" />
                <RESULT resultid="2312" eventid="70" swimtime="00:00:23.90" lane="3" heatid="70001" points="600" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100" birthdate="2017-01-01" gender="M" lastname="von Thun" firstname="Oliver" license="501090">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:58.79" heatid="4011" lane="1" />
                <ENTRY eventid="6" entrytime="00:02:09.50" heatid="6007" lane="3" />
                <ENTRY eventid="8" entrytime="00:01:03.83" heatid="8001" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:56.33" heatid="16006" lane="2" />
                <ENTRY eventid="18" entrytime="00:01:04.00" heatid="18010" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:53.55" heatid="20017" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="468" eventid="4" swimtime="00:00:50.88" lane="1" heatid="4011" points="82" />
                <RESULT resultid="469" eventid="6" swimtime="00:02:11.25" lane="3" heatid="6007" points="74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="470" eventid="8" swimtime="00:00:48.93" lane="3" heatid="8001" points="69" />
                <RESULT resultid="471" eventid="16" swimtime="00:01:53.45" lane="2" heatid="16006" points="77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="472" eventid="18" status="DSQ" swimtime="00:01:00.61" lane="3" heatid="18010" comment="Beim Anschlag an der Wende hat der Sportler nicht mit beiden Händen gleichzeitig angeschlagen." />
                <RESULT resultid="473" eventid="20" swimtime="00:01:55.57" lane="1" heatid="20017" points="58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101" birthdate="2012-01-01" gender="F" lastname="Wandschneider" firstname="Marie" license="436844">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:33.24" heatid="43005" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:47.19" heatid="27001" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:22.90" heatid="47004" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:39.69" heatid="41002" lane="2" />
                <ENTRY eventid="25" entrytime="00:00:38.53" heatid="25005" lane="4" />
                <ENTRY eventid="45" entrytime="00:01:43.26" heatid="45001" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:14.24" heatid="31005" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="474" eventid="43" swimtime="00:00:33.70" lane="1" heatid="43005" points="315" />
                <RESULT resultid="475" eventid="27" swimtime="00:00:45.53" lane="3" heatid="27001" points="241" />
                <RESULT resultid="476" eventid="47" swimtime="00:01:23.67" lane="1" heatid="47004" points="282">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="477" eventid="41" swimtime="00:00:39.89" lane="2" heatid="41002" points="228" />
                <RESULT resultid="478" eventid="25" swimtime="00:00:39.10" lane="4" heatid="25005" points="269" />
                <RESULT resultid="479" eventid="45" swimtime="00:01:42.15" lane="2" heatid="45001" points="227">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="480" eventid="31" swimtime="00:01:19.35" lane="4" heatid="31005" points="253">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102" birthdate="2017-01-01" gender="M" lastname="Wegener" firstname="Anton" license="501091">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:59.27" heatid="4011" lane="4" />
                <ENTRY eventid="6" entrytime="00:02:12.15" heatid="6007" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:48.39" heatid="8020" lane="4" />
                <ENTRY eventid="16" entrytime="00:01:57.94" heatid="16006" lane="1" />
                <ENTRY eventid="18" entrytime="00:01:06.73" heatid="18001" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:54.04" heatid="20017" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="481" eventid="4" swimtime="00:00:54.20" lane="4" heatid="4011" points="67" />
                <RESULT resultid="482" eventid="6" swimtime="00:02:22.35" lane="1" heatid="6007" points="58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="483" eventid="8" swimtime="00:00:49.17" lane="4" heatid="8020" points="68" />
                <RESULT resultid="484" eventid="16" swimtime="00:01:56.01" lane="1" heatid="16006" points="72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="485" eventid="18" swimtime="00:01:08.20" lane="2" heatid="18001" points="48" />
                <RESULT resultid="486" eventid="20" swimtime="00:01:55.99" lane="4" heatid="20017" points="57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="103" birthdate="2011-01-01" gender="F" lastname="Wilhelm" firstname="Linda" license="436850">
              <ENTRIES>
                <ENTRY eventid="29" entrytime="00:01:37.82" heatid="29004" lane="1" />
                <ENTRY eventid="47" entrytime="00:01:28.60" heatid="47005" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:27.02" heatid="33004" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:38.48" heatid="41009" lane="4" />
                <ENTRY eventid="25" entrytime="00:00:39.39" heatid="25002" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:15.24" heatid="31004" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="487" eventid="29" swimtime="00:01:30.27" lane="1" heatid="29004" points="214">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="488" eventid="47" swimtime="00:01:24.92" lane="4" heatid="47005" points="270">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="489" eventid="33" swimtime="00:01:25.99" lane="4" heatid="33004" points="283">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="490" eventid="41" swimtime="00:00:37.58" lane="4" heatid="41009" points="273" />
                <RESULT resultid="491" eventid="25" swimtime="00:00:38.68" lane="3" heatid="25002" points="278" />
                <RESULT resultid="492" eventid="31" swimtime="00:01:15.67" lane="2" heatid="31004" points="292">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:02.50" lane="3" heatid="11003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="279" eventid="11" swimtime="00:02:07.27" lane="3" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:00.67" />
                    <SPLIT distance="150" swimtime="00:01:33.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="95" number="1" />
                    <RELAYPOSITION athleteid="98" number="2" />
                    <RELAYPOSITION athleteid="71" number="3" />
                    <RELAYPOSITION athleteid="80" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="23" entrytime="00:02:22.00" lane="1" heatid="23003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="280" eventid="23" swimtime="00:02:21.75" lane="1" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:16.69" />
                    <SPLIT distance="150" swimtime="00:01:48.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="98" number="1" />
                    <RELAYPOSITION athleteid="81" number="2" />
                    <RELAYPOSITION athleteid="95" number="3" />
                    <RELAYPOSITION athleteid="71" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:01:57.00" lane="2" heatid="39003" />
                <ENTRY eventid="71" entrytime="00:02:08.50" lane="2" heatid="71003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="281" eventid="39" swimtime="00:01:57.56" lane="2" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="100" swimtime="00:00:58.27" />
                    <SPLIT distance="150" swimtime="00:01:28.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="86" number="1" />
                    <RELAYPOSITION athleteid="78" number="2" />
                    <RELAYPOSITION athleteid="91" number="3" />
                    <RELAYPOSITION athleteid="83" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="283" eventid="71" swimtime="00:02:11.24" lane="2" heatid="71003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                    <SPLIT distance="150" swimtime="00:01:41.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="86" number="1" />
                    <RELAYPOSITION athleteid="79" number="2" />
                    <RELAYPOSITION athleteid="83" number="3" />
                    <RELAYPOSITION athleteid="78" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:38.00" lane="2" heatid="40003" />
                <ENTRY eventid="72" entrytime="00:01:48.00" lane="2" heatid="72003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="282" eventid="40" swimtime="00:01:37.40" lane="2" heatid="40003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="100" swimtime="00:00:48.74" />
                    <SPLIT distance="150" swimtime="00:01:14.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="87" number="1" />
                    <RELAYPOSITION athleteid="96" number="2" />
                    <RELAYPOSITION athleteid="93" number="3" />
                    <RELAYPOSITION athleteid="99" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="284" eventid="72" swimtime="00:01:47.82" lane="2" heatid="72003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.74" />
                    <SPLIT distance="100" swimtime="00:00:57.58" />
                    <SPLIT distance="150" swimtime="00:01:23.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="99" number="1" />
                    <RELAYPOSITION athleteid="93" number="2" />
                    <RELAYPOSITION athleteid="96" number="3" />
                    <RELAYPOSITION athleteid="87" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SV Fortschritt Pirna" nation="GER" region="12" code="3387">
          <ATHLETES>
            <ATHLETE athleteid="149" birthdate="2015-01-01" gender="M" lastname="Beger" firstname="Flavius Eugen" license="492195" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:49.60" heatid="4006" lane="1" />
                <ENTRY eventid="6" entrytime="00:00:00.00" heatid="6001" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:46.91" heatid="8004" lane="3" />
                <ENTRY eventid="16" entrytime="00:00:00.00" heatid="16001" lane="1" />
                <ENTRY eventid="18" entrytime="00:01:02.35" heatid="18002" lane="1" />
                <ENTRY eventid="20" entrytime="00:00:00.00" heatid="20001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="684" eventid="4" swimtime="00:00:46.32" lane="1" heatid="4006" points="108" />
                <RESULT resultid="685" eventid="6" swimtime="00:02:14.34" lane="1" heatid="6001" points="69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="686" eventid="8" swimtime="00:00:42.70" lane="3" heatid="8004" points="105" />
                <RESULT resultid="687" eventid="16" swimtime="00:01:47.10" lane="1" heatid="16001" points="91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="688" eventid="18" status="DSQ" swimtime="00:00:56.93" lane="1" heatid="18002" comment="Der Sportler führte nach dem Start mit den Beinen wechselseitig Bewegungen aus." />
                <RESULT resultid="689" eventid="20" swimtime="00:01:43.08" lane="1" heatid="20001" points="82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150" birthdate="2017-01-01" gender="F" lastname="Haenisch" firstname="Luise" license="508206" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:01:05.76" heatid="3001" lane="3" />
                <ENTRY eventid="5" entrytime="00:00:00.00" heatid="5002" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:55.00" heatid="7003" lane="2" />
                <ENTRY eventid="15" entrytime="00:00:00.00" heatid="15003" lane="4" />
                <ENTRY eventid="17" entrytime="00:01:08.23" heatid="17003" lane="3" />
                <ENTRY eventid="19" entrytime="00:00:00.00" heatid="19001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="690" eventid="3" swimtime="00:00:59.11" lane="3" heatid="3001" points="77" />
                <RESULT resultid="691" eventid="5" status="DSQ" swimtime="00:02:15.45" lane="4" heatid="5002" comment="Beim Anschlag an der dritten Wende hat die Sportlerin nicht mit beiden Händen gleichzeitig angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="692" eventid="7" swimtime="00:00:52.99" lane="2" heatid="7003" points="81" />
                <RESULT resultid="693" eventid="15" swimtime="00:02:10.26" lane="4" heatid="15003" points="74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="694" eventid="17" swimtime="00:01:00.66" lane="3" heatid="17003" points="102" />
                <RESULT resultid="695" eventid="19" swimtime="00:01:59.88" lane="3" heatid="19001" points="73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="151" birthdate="2016-01-01" gender="F" lastname="Steiner" firstname="Frieda" license="492196" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:50.17" heatid="3009" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:46.45" heatid="7010" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:53.31" heatid="9003" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:56.61" heatid="13002" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:50.00" heatid="15006" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:44.48" heatid="19007" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="696" eventid="3" swimtime="00:00:46.04" lane="2" heatid="3009" points="164" />
                <RESULT resultid="697" eventid="7" swimtime="00:00:38.96" lane="1" heatid="7010" points="203" />
                <RESULT resultid="698" eventid="9" status="DSQ" swimtime="00:01:44.52" lane="2" heatid="9003" comment="Die Sportlerin startete vor dem Startsignal">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="699" eventid="13" swimtime="00:00:46.94" lane="1" heatid="13002" points="140" />
                <RESULT resultid="700" eventid="15" swimtime="00:01:43.72" lane="3" heatid="15006" points="148">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="701" eventid="19" swimtime="00:01:34.23" lane="3" heatid="19007" points="151">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Würzburg 05" nation="GER" region="2" code="4339">
          <ATHLETES>
            <ATHLETE athleteid="36" birthdate="2009-01-01" gender="M" lastname="Schmidt" firstname="Till Melvin" license="404171" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.61" heatid="44008" lane="1" />
                <ENTRY eventid="30" entrytime="00:01:07.29" heatid="30002" lane="3" />
                <ENTRY eventid="52" entrytime="00:02:09.78" heatid="52005" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:00.44" heatid="32007" lane="1" />
                <ENTRY eventid="50" entrytime="00:02:28.80" heatid="50002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="132" eventid="44" swimtime="00:00:27.38" lane="1" heatid="44008" points="399" />
                <RESULT resultid="133" eventid="30" swimtime="00:01:07.15" lane="3" heatid="30002" points="360">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="134" eventid="52" swimtime="00:02:09.54" lane="1" heatid="52005" points="451">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:01.89" />
                    <SPLIT distance="150" swimtime="00:01:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="135" eventid="32" swimtime="00:00:59.41" lane="1" heatid="32007" points="429">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="136" eventid="50" swimtime="00:02:26.70" lane="4" heatid="50002" points="386">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:09.50" />
                    <SPLIT distance="150" swimtime="00:01:48.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Zwickau von 1904" nation="GER" region="12" code="3400">
          <ATHLETES>
            <ATHLETE athleteid="298" birthdate="2016-01-01" gender="F" lastname="Alte" firstname="Edda Christina" license="479567" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:47.40" heatid="3011" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:42.15" heatid="7013" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:45.03" heatid="9015" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:50.93" heatid="13004" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:41.98" heatid="15016" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:39.78" heatid="19009" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1289" eventid="3" swimtime="00:00:45.93" lane="2" heatid="3011" points="166" />
                <RESULT resultid="1290" eventid="7" swimtime="00:00:40.91" lane="2" heatid="7013" points="176" />
                <RESULT resultid="1291" eventid="9" swimtime="00:01:45.01" lane="4" heatid="9015" points="155">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1292" eventid="13" swimtime="00:00:54.45" lane="4" heatid="13004" points="89" />
                <RESULT resultid="1293" eventid="15" swimtime="00:01:40.41" lane="1" heatid="15016" points="163">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1294" eventid="19" swimtime="00:01:33.49" lane="3" heatid="19009" points="155">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="299" birthdate="2017-01-01" gender="F" lastname="Bienst" firstname="Merle" license="498571">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:49.17" heatid="3019" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:51.15" heatid="7005" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:50.00" heatid="9014" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:54.30" heatid="13012" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:55.40" heatid="15015" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1295" eventid="3" swimtime="00:00:47.64" lane="3" heatid="3019" points="148" />
                <RESULT resultid="1296" eventid="7" swimtime="00:00:45.00" lane="2" heatid="7005" points="132" />
                <RESULT resultid="1297" eventid="9" swimtime="00:01:47.95" lane="1" heatid="9014" points="143">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1298" eventid="13" swimtime="00:00:54.98" lane="1" heatid="13012" points="87" />
                <RESULT resultid="1299" eventid="15" swimtime="00:01:47.85" lane="1" heatid="15015" points="131">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="300" birthdate="2015-01-01" gender="F" lastname="Birzer" firstname="Frieda" license="466284" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:33.56" heatid="5013" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:34.48" heatid="7028" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:26.24" heatid="9016" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:28.07" heatid="15017" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:43.43" heatid="17018" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:16.36" heatid="19023" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1300" eventid="5" swimtime="00:01:32.27" lane="2" heatid="5013" points="308">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1301" eventid="7" swimtime="00:00:34.09" lane="2" heatid="7028" points="304" />
                <RESULT resultid="1302" eventid="9" swimtime="00:01:25.38" lane="2" heatid="9016" points="289">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1303" eventid="15" swimtime="00:01:24.83" lane="1" heatid="15017" points="270">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1304" eventid="17" swimtime="00:00:43.11" lane="2" heatid="17018" points="284" />
                <RESULT resultid="1305" eventid="19" swimtime="00:01:15.25" lane="2" heatid="19023" points="297">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="301" birthdate="2013-01-01" gender="F" lastname="Dressel" firstname="Clara" license="447504" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:35.70" heatid="5015" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:34.66" heatid="7025" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:26.05" heatid="15019" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:43.67" heatid="17020" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1306" eventid="5" swimtime="00:01:33.46" lane="4" heatid="5015" points="297">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1307" eventid="7" swimtime="00:00:34.43" lane="4" heatid="7025" points="295" />
                <RESULT resultid="1308" eventid="15" swimtime="00:01:24.86" lane="4" heatid="15019" points="270">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1309" eventid="17" swimtime="00:00:44.07" lane="1" heatid="17020" points="266" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="302" birthdate="2017-01-01" gender="M" lastname="Dressel" firstname="Johann" license="496421">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:02:05.00" heatid="6007" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:54.38" heatid="8002" lane="3" />
                <ENTRY eventid="10" entrytime="00:02:00.00" heatid="10008" lane="2" />
                <ENTRY eventid="18" entrytime="00:01:04.84" heatid="18010" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:55.00" heatid="20002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1310" eventid="6" swimtime="00:02:10.27" lane="2" heatid="6007" points="76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1311" eventid="8" swimtime="00:00:50.10" lane="3" heatid="8002" points="65" />
                <RESULT resultid="1312" eventid="10" swimtime="00:02:05.62" lane="2" heatid="10008" points="60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1313" eventid="18" swimtime="00:01:01.25" lane="4" heatid="18010" points="67" />
                <RESULT resultid="1314" eventid="20" swimtime="00:01:58.95" lane="3" heatid="20002" points="53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="303" birthdate="2015-01-01" gender="F" lastname="Dusl" firstname="Mara" license="466278" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.45" heatid="3015" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:40.80" heatid="7015" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:41.43" heatid="9006" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:34.79" heatid="15012" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:55.34" heatid="17006" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:32.37" heatid="19012" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1315" eventid="3" swimtime="00:00:45.37" lane="4" heatid="3015" points="172" />
                <RESULT resultid="1316" eventid="7" swimtime="00:00:40.51" lane="4" heatid="7015" points="181" />
                <RESULT resultid="1317" eventid="9" swimtime="00:01:39.73" lane="1" heatid="9006" points="181">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1318" eventid="15" swimtime="00:01:38.78" lane="4" heatid="15012" points="171">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1319" eventid="17" swimtime="00:00:55.14" lane="3" heatid="17006" points="136" />
                <RESULT resultid="1320" eventid="19" swimtime="00:01:34.27" lane="3" heatid="19012" points="151">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="304" birthdate="2013-01-01" gender="F" lastname="Fenzel" firstname="Valeria" license="448580" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:32.00" heatid="1005" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:34.11" heatid="7030" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:25.49" heatid="9013" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:39.73" heatid="13011" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:26.34" heatid="15014" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:14.22" heatid="19025" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1321" eventid="1" swimtime="00:01:31.16" lane="3" heatid="1005" points="208">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1322" eventid="7" swimtime="00:00:33.27" lane="4" heatid="7030" points="327" />
                <RESULT resultid="1323" eventid="9" swimtime="00:01:25.97" lane="2" heatid="9013" points="284">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1324" eventid="13" swimtime="00:00:39.28" lane="1" heatid="13011" points="239" />
                <RESULT resultid="1325" eventid="15" swimtime="00:01:26.22" lane="4" heatid="15014" points="258">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1326" eventid="19" swimtime="00:01:14.66" lane="1" heatid="19025" points="304">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="305" birthdate="2008-01-01" gender="M" lastname="Filiz" firstname="Denis" license="363786" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.37" heatid="44009" lane="2" />
                <ENTRY eventid="48" entrytime="00:01:08.54" heatid="48005" lane="4" />
                <ENTRY eventid="34" entrytime="00:01:09.75" heatid="34008" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:30.24" heatid="26005" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1327" eventid="44" swimtime="00:00:27.13" lane="2" heatid="44009" points="410" />
                <RESULT resultid="1328" eventid="48" swimtime="00:01:09.00" lane="4" heatid="48005" points="343">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1329" eventid="34" swimtime="00:01:10.27" lane="3" heatid="34008" points="344">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1330" eventid="26" swimtime="00:00:30.86" lane="4" heatid="26005" points="367" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="306" birthdate="2014-01-01" gender="F" lastname="Fischer" firstname="Alma" license="461986" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:48.10" heatid="5006" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:44.22" heatid="7011" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:38.47" heatid="9007" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:51.04" heatid="13003" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:49.82" heatid="17011" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:31.75" heatid="19013" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1331" eventid="5" swimtime="00:01:43.47" lane="2" heatid="5006" points="218">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1332" eventid="7" swimtime="00:00:39.20" lane="1" heatid="7011" points="200" />
                <RESULT resultid="1333" eventid="9" swimtime="00:01:37.69" lane="4" heatid="9007" points="193">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1334" eventid="13" swimtime="00:00:46.29" lane="2" heatid="13003" points="146" />
                <RESULT resultid="1335" eventid="17" swimtime="00:00:48.30" lane="4" heatid="17011" points="202" />
                <RESULT resultid="1336" eventid="19" swimtime="00:01:31.47" lane="4" heatid="19013" points="165">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="307" birthdate="2017-01-01" gender="F" lastname="Frank" firstname="Lorelei" license="498012">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:52.79" heatid="5011" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:48.39" heatid="7008" lane="1" />
                <ENTRY eventid="9" entrytime="00:02:00.00" heatid="9003" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:50.00" heatid="13012" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:53.30" heatid="17016" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:50.27" heatid="19005" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1337" eventid="5" swimtime="00:01:47.10" lane="2" heatid="5011" points="197">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1338" eventid="7" swimtime="00:00:50.29" lane="1" heatid="7008" points="94" />
                <RESULT resultid="1339" eventid="9" swimtime="00:01:46.86" lane="4" heatid="9003" points="147">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1340" eventid="13" swimtime="00:00:55.33" lane="3" heatid="13012" points="85" />
                <RESULT resultid="1341" eventid="17" swimtime="00:00:52.36" lane="3" heatid="17016" points="159" />
                <RESULT resultid="1342" eventid="19" swimtime="00:01:47.63" lane="4" heatid="19005" points="101">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="308" birthdate="1990-01-01" gender="M" lastname="Hahn" firstname="Renè" license="139403">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:25.57" heatid="44012" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:33.56" heatid="28006" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:27.91" heatid="42008" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1343" eventid="44" swimtime="00:00:25.03" lane="3" heatid="44012" points="522" />
                <RESULT resultid="1344" eventid="28" swimtime="00:00:34.15" lane="3" heatid="28006" points="389" />
                <RESULT resultid="1345" eventid="42" swimtime="00:00:27.88" lane="4" heatid="42008" points="474" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="309" birthdate="2010-01-01" gender="M" lastname="Käser" firstname="Mika Marco" license="423052" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:28.95" heatid="44006" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:37.72" heatid="28004" lane="3" />
                <ENTRY eventid="52" entrytime="00:02:24.83" heatid="52004" lane="4" />
                <ENTRY eventid="38" entrytime="00:03:07.00" heatid="38004" lane="4" />
                <ENTRY eventid="32" entrytime="00:01:04.18" heatid="32005" lane="4" />
                <ENTRY eventid="54" entrytime="00:02:48.41" heatid="54002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1346" eventid="44" swimtime="00:00:27.93" lane="1" heatid="44006" points="376" />
                <RESULT resultid="1347" eventid="28" swimtime="00:00:37.61" lane="3" heatid="28004" points="291" />
                <RESULT resultid="1348" eventid="52" swimtime="00:02:24.09" lane="4" heatid="52004" points="327">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1349" eventid="38" swimtime="00:02:59.43" lane="4" heatid="38004" points="300">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                    <SPLIT distance="100" swimtime="00:01:26.06" />
                    <SPLIT distance="150" swimtime="00:02:12.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1350" eventid="32" swimtime="00:01:05.08" lane="4" heatid="32005" points="327">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1351" eventid="54" swimtime="00:02:44.03" lane="3" heatid="54002" points="298">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:02:08.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="310" birthdate="2012-01-01" gender="F" lastname="Komar" firstname="Lindsay" license="436924" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.22" heatid="43010" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:40.31" heatid="27006" lane="3" />
                <ENTRY eventid="29" entrytime="00:01:17.84" heatid="29003" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:16.42" heatid="33006" lane="2" />
                <ENTRY eventid="67" entrytime="00:00:29.46" heatid="67000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1352" eventid="43" swimtime="00:00:29.46" lane="3" heatid="43010" points="471" />
                <RESULT resultid="1353" eventid="27" swimtime="00:00:39.41" lane="3" heatid="27006" points="373" />
                <RESULT resultid="1354" eventid="29" swimtime="00:01:18.74" lane="3" heatid="29003" points="323">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1355" eventid="33" swimtime="00:01:16.90" lane="2" heatid="33006" points="396">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2298" eventid="67" status="WDR" swimtime="00:00:00.00" lane="0" heatid="67000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="311" birthdate="2007-01-01" gender="F" lastname="Kunz" firstname="Jenny" license="363787" nation="GER">
              <ENTRIES>
                <ENTRY eventid="29" entrytime="00:01:13.80" heatid="29006" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:17.05" heatid="47007" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:09.49" heatid="31006" lane="2" />
                <ENTRY eventid="35" entrytime="00:02:44.14" heatid="35003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1356" eventid="29" swimtime="00:01:15.93" lane="3" heatid="29006" points="360">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1357" eventid="47" swimtime="00:01:17.07" lane="3" heatid="47007" points="361">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1358" eventid="31" swimtime="00:01:09.30" lane="2" heatid="31006" points="381">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1359" eventid="35" swimtime="00:02:49.35" lane="1" heatid="35003" points="346">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:21.01" />
                    <SPLIT distance="150" swimtime="00:02:06.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="312" birthdate="2005-01-01" gender="M" lastname="Kunz" firstname="Jeremy" license="348770" nation="GER">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:31.29" heatid="28011" lane="1" />
                <ENTRY eventid="30" entrytime="00:00:57.67" heatid="30006" lane="3" />
                <ENTRY eventid="34" entrytime="00:00:58.78" heatid="34009" lane="1" />
                <ENTRY eventid="52" entrytime="00:01:52.82" heatid="52006" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:26.78" heatid="42009" lane="1" />
                <ENTRY eventid="26" entrytime="00:00:27.02" heatid="26010" lane="4" />
                <ENTRY eventid="32" entrytime="00:00:52.92" heatid="32013" lane="1" />
                <ENTRY eventid="36" entrytime="00:02:04.14" heatid="36003" lane="2" />
                <ENTRY eventid="54" entrytime="00:02:08.60" heatid="54005" lane="3" />
                <ENTRY eventid="62" entrytime="00:00:30.60" heatid="62001" lane="4" />
                <ENTRY eventid="58" entrytime="00:00:27.24" heatid="58001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1360" eventid="28" swimtime="00:00:30.60" lane="1" heatid="28011" points="542" />
                <RESULT resultid="1361" eventid="30" swimtime="00:00:58.27" lane="3" heatid="30006" points="551">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1362" eventid="34" swimtime="00:00:59.19" lane="1" heatid="34009" points="577">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1363" eventid="52" swimtime="00:02:00.96" lane="2" heatid="52006" points="554">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                    <SPLIT distance="100" swimtime="00:00:58.98" />
                    <SPLIT distance="150" swimtime="00:01:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1364" eventid="42" swimtime="00:00:26.81" lane="1" heatid="42009" points="533" />
                <RESULT resultid="1365" eventid="26" swimtime="00:00:27.24" lane="4" heatid="26010" points="534" />
                <RESULT resultid="1366" eventid="32" swimtime="00:00:53.89" lane="1" heatid="32013" points="576">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1367" eventid="36" swimtime="00:02:18.84" lane="2" heatid="36003" points="440">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:08.75" />
                    <SPLIT distance="150" swimtime="00:01:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1368" eventid="54" swimtime="00:02:18.44" lane="3" heatid="54005" points="496">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="100" swimtime="00:01:05.29" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2362" eventid="58" swimtime="00:00:27.18" lane="4" heatid="58001" points="538" />
                <RESULT resultid="2330" eventid="62" swimtime="00:00:30.88" lane="4" heatid="62001" points="527" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="313" birthdate="2017-01-01" gender="F" lastname="Landgraf" firstname="Emma" license="496724">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:01:00.58" heatid="3002" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:57.54" heatid="7003" lane="4" />
                <ENTRY eventid="9" entrytime="00:02:00.00" heatid="9002" lane="2" />
                <ENTRY eventid="13" entrytime="00:01:01.43" heatid="13001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1369" eventid="3" swimtime="00:00:54.75" lane="1" heatid="3002" points="98" />
                <RESULT resultid="1370" eventid="7" swimtime="00:00:53.41" lane="4" heatid="7003" points="79" />
                <RESULT resultid="1371" eventid="9" swimtime="00:02:01.68" lane="2" heatid="9002" points="100">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1372" eventid="13" swimtime="00:01:03.17" lane="2" heatid="13001" points="57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="314" birthdate="2015-01-01" gender="F" lastname="Lemke" firstname="Lilly-Rose" license="466280" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:45.21" heatid="3014" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:41.25" heatid="7014" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:39.30" heatid="9006" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:40.85" heatid="15009" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:54.78" heatid="17007" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:34.65" heatid="19011" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1373" eventid="3" swimtime="00:00:42.99" lane="1" heatid="3014" points="202" />
                <RESULT resultid="1374" eventid="7" swimtime="00:00:38.49" lane="3" heatid="7014" points="211" />
                <RESULT resultid="1375" eventid="9" swimtime="00:01:41.78" lane="3" heatid="9006" points="171">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1376" eventid="15" swimtime="00:01:36.99" lane="4" heatid="15009" points="181">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1377" eventid="17" swimtime="00:00:53.85" lane="4" heatid="17007" points="146" />
                <RESULT resultid="1378" eventid="19" swimtime="00:01:34.94" lane="1" heatid="19011" points="148">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="315" birthdate="2009-01-01" gender="F" lastname="Nahlovsky" firstname="Lilly" license="410485" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:28.42" heatid="43012" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:36.90" heatid="27005" lane="2" />
                <ENTRY eventid="47" entrytime="00:01:10.77" heatid="47006" lane="1" />
                <ENTRY eventid="33" entrytime="00:01:12.34" heatid="33008" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:31.31" heatid="41007" lane="2" />
                <ENTRY eventid="25" entrytime="00:00:31.38" heatid="25007" lane="3" />
                <ENTRY eventid="68" entrytime="00:00:28.26" heatid="68001" lane="4" />
                <ENTRY eventid="59" entrytime="00:00:36.72" heatid="59001" lane="2" />
                <ENTRY eventid="64" entrytime="00:00:31.13" heatid="64001" lane="4" />
                <ENTRY eventid="56" entrytime="00:00:31.84" heatid="56001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1379" eventid="43" swimtime="00:00:28.26" lane="4" heatid="43012" points="534" />
                <RESULT resultid="1380" eventid="27" swimtime="00:00:36.72" lane="2" heatid="27005" points="461" />
                <RESULT resultid="1381" eventid="47" swimtime="00:01:10.05" lane="1" heatid="47006" points="481">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1382" eventid="33" swimtime="00:01:12.76" lane="1" heatid="33008" points="468">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1383" eventid="41" swimtime="00:00:31.13" lane="2" heatid="41007" points="480" />
                <RESULT resultid="1384" eventid="25" swimtime="00:00:31.84" lane="3" heatid="25007" points="498" />
                <RESULT resultid="2352" eventid="56" swimtime="00:00:31.31" lane="3" heatid="56001" points="524" />
                <RESULT resultid="2315" eventid="59" swimtime="00:00:36.42" lane="2" heatid="59001" points="472" />
                <RESULT resultid="2338" eventid="64" swimtime="00:00:30.97" lane="4" heatid="64001" points="487" />
                <RESULT resultid="2306" eventid="68" swimtime="00:00:28.38" lane="4" heatid="68001" points="527" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="316" birthdate="2013-01-01" gender="F" lastname="Navarro Perez" firstname="Angielina" license="494142" nation="ESP">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:43.05" heatid="3016" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:37.06" heatid="7019" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:30.77" heatid="9011" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:40.52" heatid="13011" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:35.62" heatid="15011" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:23.81" heatid="19016" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1385" eventid="3" swimtime="00:00:41.37" lane="2" heatid="3016" points="227" />
                <RESULT resultid="1386" eventid="7" swimtime="00:00:36.89" lane="2" heatid="7019" points="240" />
                <RESULT resultid="1387" eventid="9" swimtime="00:01:31.41" lane="2" heatid="9011" points="236">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1388" eventid="13" swimtime="00:00:42.04" lane="4" heatid="13011" points="195" />
                <RESULT resultid="1389" eventid="15" swimtime="00:01:34.35" lane="2" heatid="15011" points="196">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1390" eventid="19" swimtime="00:01:23.62" lane="3" heatid="19016" points="217">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="317" birthdate="2015-01-01" gender="F" lastname="Navarro Perez" firstname="Arianna" license="494141" nation="ESP">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:50.00" heatid="1001" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:43.24" heatid="7012" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:45.80" heatid="9004" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:48.21" heatid="13005" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:43.61" heatid="15008" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:36.34" heatid="19010" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1391" eventid="1" swimtime="00:01:53.07" lane="3" heatid="1001" points="109">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1392" eventid="7" swimtime="00:00:42.33" lane="4" heatid="7012" points="158" />
                <RESULT resultid="1393" eventid="9" swimtime="00:01:41.10" lane="3" heatid="9004" points="174">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1394" eventid="13" swimtime="00:00:48.73" lane="3" heatid="13005" points="125" />
                <RESULT resultid="1395" eventid="15" swimtime="00:01:42.50" lane="3" heatid="15008" points="153">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1396" eventid="19" swimtime="00:01:34.31" lane="3" heatid="19010" points="151">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="318" birthdate="2012-01-01" gender="M" lastname="Nawrath" firstname="Jonas" license="443627" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:26.94" heatid="6012" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:30.44" heatid="8025" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:18.80" heatid="10013" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:31.30" heatid="14012" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:37.33" heatid="18015" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:09.75" heatid="20016" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1397" eventid="6" swimtime="00:01:24.33" lane="4" heatid="6012" points="281">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1398" eventid="8" swimtime="00:00:28.97" lane="1" heatid="8025" points="336" />
                <RESULT resultid="1399" eventid="10" swimtime="00:01:17.24" lane="1" heatid="10013" points="259">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1400" eventid="14" swimtime="00:00:31.27" lane="3" heatid="14012" points="336" />
                <RESULT resultid="1401" eventid="18" swimtime="00:00:36.26" lane="3" heatid="18015" points="325" />
                <RESULT resultid="1402" eventid="20" swimtime="00:01:09.78" lane="2" heatid="20016" points="265">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="319" birthdate="2017-01-01" gender="F" lastname="Oehler" firstname="Magdalena" license="496426">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:57.00" heatid="3000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:52.06" heatid="7000" lane="0" />
                <ENTRY eventid="9" entrytime="00:02:00.00" heatid="9000" lane="0" />
                <ENTRY eventid="13" entrytime="00:01:00.50" heatid="13000" lane="0" />
                <ENTRY eventid="17" entrytime="00:00:57.00" heatid="17000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1403" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="1404" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="1405" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
                <RESULT resultid="1406" eventid="13" status="WDR" swimtime="00:00:00.00" lane="0" heatid="13000" />
                <RESULT resultid="1407" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="320" birthdate="2014-01-01" gender="F" lastname="Paul" firstname="Ilvy" license="464150" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:32.60" heatid="1002" lane="3" />
                <ENTRY eventid="5" entrytime="00:01:33.05" heatid="5014" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:26.33" heatid="9013" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:36.35" heatid="13015" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:42.20" heatid="17019" lane="2" />
                <ENTRY eventid="21" entrytime="00:03:12.57" heatid="21003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1408" eventid="1" swimtime="00:01:31.19" lane="3" heatid="1002" points="208">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1409" eventid="5" swimtime="00:01:31.66" lane="3" heatid="5014" points="314">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1410" eventid="9" swimtime="00:01:23.71" lane="3" heatid="9013" points="307">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1411" eventid="13" swimtime="00:00:38.33" lane="1" heatid="13015" points="257" />
                <RESULT resultid="1412" eventid="17" swimtime="00:00:39.17" lane="2" heatid="17019" points="379" />
                <RESULT resultid="1413" eventid="21" swimtime="00:03:09.46" lane="3" heatid="21003" points="266">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:30.17" />
                    <SPLIT distance="150" swimtime="00:02:24.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="321" birthdate="2004-01-01" gender="M" lastname="Paul" firstname="Lenny" license="331135" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:25.84" heatid="44012" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:32.43" heatid="28007" lane="3" />
                <ENTRY eventid="30" entrytime="00:01:02.42" heatid="30003" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:26.90" heatid="42009" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:30.19" heatid="26005" lane="1" />
                <ENTRY eventid="32" entrytime="00:00:58.17" heatid="32009" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1414" eventid="44" swimtime="00:00:26.62" lane="1" heatid="44012" points="434" />
                <RESULT resultid="1415" eventid="28" swimtime="00:00:33.30" lane="3" heatid="28007" points="420" />
                <RESULT resultid="1416" eventid="30" swimtime="00:01:03.45" lane="3" heatid="30003" points="427">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1417" eventid="42" swimtime="00:00:28.01" lane="4" heatid="42009" points="468" />
                <RESULT resultid="1418" eventid="26" swimtime="00:00:30.84" lane="1" heatid="26005" points="368" />
                <RESULT resultid="1419" eventid="32" swimtime="00:01:01.58" lane="1" heatid="32009" points="386">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="322" birthdate="2014-01-01" gender="M" lastname="Plettig" firstname="Ben" license="464151" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:28.02" heatid="2002" lane="2" />
                <ENTRY eventid="4" entrytime="00:00:36.55" heatid="4014" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:33.81" heatid="8017" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:38.26" heatid="14006" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:19.11" heatid="16009" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:13.16" heatid="20016" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1420" eventid="2" swimtime="00:01:26.84" lane="2" heatid="2002" points="166">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1421" eventid="4" swimtime="00:00:35.52" lane="2" heatid="4014" points="241" />
                <RESULT resultid="1422" eventid="8" swimtime="00:00:33.31" lane="3" heatid="8017" points="221" />
                <RESULT resultid="1423" eventid="14" swimtime="00:00:36.50" lane="3" heatid="14006" points="211" />
                <RESULT resultid="1424" eventid="16" swimtime="00:01:19.31" lane="2" heatid="16009" points="226">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1425" eventid="20" swimtime="00:01:14.11" lane="4" heatid="20016" points="221">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="323" birthdate="2016-01-01" gender="F" lastname="Plettig" firstname="Lena" license="479565" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:48.14" heatid="3010" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:38.95" heatid="7018" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:42.03" heatid="9015" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:43.06" heatid="13013" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:52.42" heatid="17009" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:33.69" heatid="19012" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1426" eventid="3" swimtime="00:00:46.18" lane="3" heatid="3010" points="163" />
                <RESULT resultid="1427" eventid="7" swimtime="00:00:40.40" lane="4" heatid="7018" points="182" />
                <RESULT resultid="1428" eventid="9" swimtime="00:01:37.15" lane="1" heatid="9015" points="196">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1429" eventid="13" swimtime="00:00:43.64" lane="1" heatid="13013" points="174" />
                <RESULT resultid="1430" eventid="17" swimtime="00:00:53.81" lane="3" heatid="17009" points="146" />
                <RESULT resultid="1431" eventid="19" swimtime="00:01:36.12" lane="4" heatid="19012" points="142">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="324" birthdate="2014-01-01" gender="F" lastname="Pöhler" firstname="Edda" license="479562" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:45.54" heatid="5007" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:39.21" heatid="7017" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:44.98" heatid="9005" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:45.98" heatid="13007" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:48.17" heatid="17012" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:31.93" heatid="19012" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1432" eventid="5" swimtime="00:01:43.47" lane="3" heatid="5007" points="218">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1433" eventid="7" swimtime="00:00:38.31" lane="1" heatid="7017" points="214" />
                <RESULT resultid="1434" eventid="9" swimtime="00:01:36.90" lane="1" heatid="9005" points="198">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1435" eventid="13" swimtime="00:00:42.65" lane="1" heatid="13007" points="186" />
                <RESULT resultid="1436" eventid="17" swimtime="00:00:47.14" lane="3" heatid="17012" points="217" />
                <RESULT resultid="1437" eventid="19" swimtime="00:01:29.15" lane="2" heatid="19012" points="179">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="325" birthdate="2013-01-01" gender="M" lastname="Richter" firstname="Luke" license="446150" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:37.27" heatid="4015" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:32.20" heatid="8019" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:21.70" heatid="10012" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:36.79" heatid="14011" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:12.58" heatid="20021" lane="4" />
                <ENTRY eventid="22" entrytime="00:02:51.22" heatid="22005" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1438" eventid="4" swimtime="00:00:36.89" lane="2" heatid="4015" points="215" />
                <RESULT resultid="1439" eventid="8" swimtime="00:00:31.69" lane="1" heatid="8019" points="257" />
                <RESULT resultid="1440" eventid="10" swimtime="00:01:20.22" lane="3" heatid="10012" points="231">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1441" eventid="14" swimtime="00:00:38.84" lane="4" heatid="14011" points="175" />
                <RESULT resultid="1442" eventid="20" swimtime="00:01:09.76" lane="4" heatid="20021" points="265">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1443" eventid="22" swimtime="00:02:58.42" lane="4" heatid="22005" points="231">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                    <SPLIT distance="100" swimtime="00:01:24.01" />
                    <SPLIT distance="150" swimtime="00:02:18.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="326" birthdate="2016-01-01" gender="F" lastname="Rödel" firstname="Anna Karla" license="499253" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:51.83" heatid="3009" lane="1" />
                <ENTRY eventid="5" entrytime="00:01:57.44" heatid="5004" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:48.61" heatid="7008" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:47.32" heatid="15007" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:54.39" heatid="17007" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:45.00" heatid="19006" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1444" eventid="3" swimtime="00:00:50.34" lane="1" heatid="3009" points="126" />
                <RESULT resultid="1445" eventid="5" swimtime="00:01:57.78" lane="1" heatid="5004" points="148">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1446" eventid="7" swimtime="00:00:46.68" lane="4" heatid="7008" points="118" />
                <RESULT resultid="1447" eventid="15" status="DSQ" swimtime="00:01:49.90" lane="4" heatid="15007" comment="Bei der zweiten Wende wurde die Wand nicht berührt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1448" eventid="17" swimtime="00:00:53.50" lane="1" heatid="17007" points="149" />
                <RESULT resultid="1449" eventid="19" swimtime="00:01:43.83" lane="1" heatid="19006" points="113">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="327" birthdate="2010-01-01" gender="F" lastname="Rohatzsch" firstname="Maxime" license="410491" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.78" heatid="43007" lane="1" />
                <ENTRY eventid="47" entrytime="00:01:16.20" heatid="47003" lane="3" />
                <ENTRY eventid="51" entrytime="00:02:36.24" heatid="51002" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:33.85" heatid="41006" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:09.45" heatid="31007" lane="4" />
                <ENTRY eventid="35" entrytime="00:02:45.70" heatid="35002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1450" eventid="43" swimtime="00:00:30.88" lane="1" heatid="43007" points="409" />
                <RESULT resultid="1451" eventid="47" swimtime="00:01:16.44" lane="3" heatid="47003" points="370">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1452" eventid="51" swimtime="00:02:30.68" lane="4" heatid="51002" points="392">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:11.09" />
                    <SPLIT distance="150" swimtime="00:01:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1453" eventid="41" swimtime="00:00:34.01" lane="4" heatid="41006" points="368" />
                <RESULT resultid="1454" eventid="31" swimtime="00:01:08.68" lane="4" heatid="31007" points="391">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1455" eventid="35" swimtime="00:02:48.29" lane="3" heatid="35002" points="353">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:02:05.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="328" birthdate="1997-01-01" gender="M" lastname="Rohmberger" firstname="Thomas" license="210024" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:23.00" heatid="44017" lane="3" />
                <ENTRY eventid="34" entrytime="00:00:55.00" heatid="34009" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:25.00" heatid="42013" lane="3" />
                <ENTRY eventid="32" entrytime="00:00:51.00" heatid="32013" lane="2" />
                <ENTRY eventid="70" entrytime="00:00:23.96" heatid="70001" lane="4" />
                <ENTRY eventid="66" entrytime="00:00:25.03" heatid="66001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1456" eventid="44" swimtime="00:00:23.96" lane="3" heatid="44017" points="595" />
                <RESULT resultid="1457" eventid="34" swimtime="00:00:59.24" lane="2" heatid="34009" points="575">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1458" eventid="42" swimtime="00:00:25.03" lane="3" heatid="42013" points="656" />
                <RESULT resultid="1459" eventid="32" swimtime="00:00:54.07" lane="2" heatid="32013" points="570">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2344" eventid="66" swimtime="00:00:24.53" lane="3" heatid="66001" points="697" />
                <RESULT resultid="2314" eventid="70" swimtime="00:00:23.85" lane="4" heatid="70001" points="603" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="329" birthdate="2015-01-01" gender="F" lastname="Rudolph" firstname="Frieda" license="471935" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:55.00" heatid="5005" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:42.67" heatid="7013" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:50.00" heatid="9004" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:49.85" heatid="13004" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:52.46" heatid="17009" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:40.00" heatid="19009" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1460" eventid="5" swimtime="00:01:53.08" lane="1" heatid="5005" points="167">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1461" eventid="7" swimtime="00:00:43.11" lane="1" heatid="7013" points="150" />
                <RESULT resultid="1462" eventid="9" swimtime="00:01:52.12" lane="4" heatid="9004" points="128">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1463" eventid="13" swimtime="00:00:48.72" lane="2" heatid="13004" points="125" />
                <RESULT resultid="1464" eventid="17" swimtime="00:00:54.06" lane="1" heatid="17009" points="144" />
                <RESULT resultid="1465" eventid="19" swimtime="00:01:43.56" lane="1" heatid="19009" points="114">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="330" birthdate="2013-01-01" gender="F" lastname="Schlawitz" firstname="Amalia" license="464149" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:41.37" heatid="3017" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:34.67" heatid="7024" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:34.38" heatid="9010" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:30.28" heatid="15012" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:16.01" heatid="19025" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1466" eventid="3" swimtime="00:00:40.36" lane="2" heatid="3017" points="244" />
                <RESULT resultid="1467" eventid="7" swimtime="00:00:34.12" lane="2" heatid="7024" points="303" />
                <RESULT resultid="1468" eventid="9" swimtime="00:01:29.45" lane="2" heatid="9010" points="252">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1469" eventid="15" swimtime="00:01:29.03" lane="2" heatid="15012" points="234">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1470" eventid="19" swimtime="00:01:14.76" lane="4" heatid="19025" points="303">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="331" birthdate="1999-01-01" gender="M" lastname="Schneider" firstname="Eric" license="242941" nation="GER">
              <ENTRIES>
                <ENTRY eventid="34" entrytime="00:01:00.44" heatid="34009" lane="4" />
                <ENTRY eventid="38" entrytime="00:02:36.33" heatid="38006" lane="4" />
                <ENTRY eventid="26" entrytime="00:00:27.73" heatid="26006" lane="2" />
                <ENTRY eventid="46" entrytime="00:01:07.86" heatid="46007" lane="3" />
                <ENTRY eventid="36" entrytime="00:02:24.60" heatid="36002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1471" eventid="34" swimtime="00:01:01.24" lane="4" heatid="34009" points="521">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1472" eventid="38" swimtime="00:02:32.78" lane="4" heatid="38006" points="486">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:12.19" />
                    <SPLIT distance="150" swimtime="00:01:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1473" eventid="26" swimtime="00:00:28.33" lane="2" heatid="26006" points="475" />
                <RESULT resultid="1474" eventid="46" swimtime="00:01:09.48" lane="3" heatid="46007" points="503">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1475" eventid="36" status="DNS" swimtime="00:00:00.00" lane="2" heatid="36002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="332" birthdate="2013-01-01" gender="F" lastname="Schneider" firstname="Laura" license="447503" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:18.35" heatid="1005" lane="2" />
                <ENTRY eventid="5" entrytime="00:01:17.71" heatid="5015" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:15.20" heatid="9018" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:33.38" heatid="13016" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:35.43" heatid="17020" lane="2" />
                <ENTRY eventid="21" entrytime="00:02:46.52" heatid="21004" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1476" eventid="1" swimtime="00:01:16.65" lane="2" heatid="1005" points="350">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1477" eventid="5" swimtime="00:01:17.50" lane="2" heatid="5015" points="520">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1478" eventid="9" swimtime="00:01:13.35" lane="2" heatid="9018" points="457">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1479" eventid="13" swimtime="00:00:32.21" lane="2" heatid="13016" points="433" />
                <RESULT resultid="1480" eventid="17" swimtime="00:00:34.98" lane="2" heatid="17020" points="533" />
                <RESULT resultid="1481" eventid="21" swimtime="00:02:45.24" lane="2" heatid="21004" points="401">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:19.28" />
                    <SPLIT distance="150" swimtime="00:02:05.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="333" birthdate="2015-01-01" gender="F" lastname="Schneider" firstname="Linda" license="466281" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:25.00" heatid="1003" lane="2" />
                <ENTRY eventid="3" entrytime="00:00:42.65" heatid="3021" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:36.19" heatid="7022" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:41.85" heatid="13014" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:32.18" heatid="15012" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:22.88" heatid="19017" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1482" eventid="1" swimtime="00:01:39.79" lane="2" heatid="1003" points="158">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1483" eventid="3" swimtime="00:00:41.60" lane="4" heatid="3021" points="223" />
                <RESULT resultid="1484" eventid="7" swimtime="00:00:35.31" lane="1" heatid="7022" points="273" />
                <RESULT resultid="1485" eventid="13" swimtime="00:00:40.43" lane="1" heatid="13014" points="219" />
                <RESULT resultid="1486" eventid="15" swimtime="00:01:31.37" lane="3" heatid="15012" points="216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1487" eventid="19" swimtime="00:01:20.78" lane="2" heatid="19017" points="240">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="334" birthdate="2014-01-01" gender="F" lastname="Sprenger" firstname="Lara" license="456271" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:38.21" heatid="3022" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:33.68" heatid="7025" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:27.07" heatid="9013" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:41.22" heatid="13010" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:20.60" heatid="15018" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:14.05" heatid="19024" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1488" eventid="3" swimtime="00:00:37.17" lane="1" heatid="3022" points="313" />
                <RESULT resultid="1489" eventid="7" swimtime="00:00:33.96" lane="2" heatid="7025" points="307" />
                <RESULT resultid="1490" eventid="9" swimtime="00:01:26.62" lane="1" heatid="9013" points="277">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1491" eventid="13" swimtime="00:00:41.65" lane="1" heatid="13010" points="200" />
                <RESULT resultid="1492" eventid="15" swimtime="00:01:21.94" lane="1" heatid="15018" points="300">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1493" eventid="19" swimtime="00:01:13.37" lane="4" heatid="19024" points="321">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="335" birthdate="2017-01-01" gender="F" lastname="Strangfeld" firstname="Ida" license="496430">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:50.67" heatid="3019" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:43.38" heatid="7026" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:49.54" heatid="9014" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:50.00" heatid="13012" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:51.99" heatid="15015" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:39.41" heatid="19021" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1494" eventid="3" swimtime="00:00:48.26" lane="4" heatid="3019" points="143" />
                <RESULT resultid="1495" eventid="7" swimtime="00:00:44.42" lane="3" heatid="7026" points="137" />
                <RESULT resultid="1496" eventid="9" swimtime="00:01:45.13" lane="3" heatid="9014" points="155">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1497" eventid="13" swimtime="00:00:54.71" lane="2" heatid="13012" points="88" />
                <RESULT resultid="1498" eventid="15" swimtime="00:01:47.37" lane="3" heatid="15015" points="133">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1499" eventid="19" status="DSQ" swimtime="00:01:39.75" lane="3" heatid="19021" comment="Die Sportlerin startete vor dem Startsignal">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="336" birthdate="2011-01-01" gender="M" lastname="Suhr" firstname="Damian" license="438666" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:29.98" heatid="44005" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:41.11" heatid="28003" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:17.67" heatid="34004" lane="4" />
                <ENTRY eventid="38" entrytime="00:03:13.00" heatid="38003" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:34.46" heatid="26007" lane="3" />
                <ENTRY eventid="32" entrytime="00:01:08.80" heatid="32004" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1500" eventid="44" swimtime="00:00:29.88" lane="4" heatid="44005" points="307" />
                <RESULT resultid="1501" eventid="28" swimtime="00:00:41.11" lane="1" heatid="28003" points="223" />
                <RESULT resultid="1502" eventid="34" swimtime="00:01:16.60" lane="4" heatid="34004" points="266">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1503" eventid="38" swimtime="00:03:12.59" lane="3" heatid="38003" points="242">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                    <SPLIT distance="100" swimtime="00:01:31.66" />
                    <SPLIT distance="150" swimtime="00:02:22.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1504" eventid="26" swimtime="00:00:33.41" lane="3" heatid="26007" points="289" />
                <RESULT resultid="1505" eventid="32" swimtime="00:01:08.23" lane="1" heatid="32004" points="283">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="337" birthdate="2004-01-01" gender="F" lastname="Süppel" firstname="Laura" license="329276" nation="GER">
              <ENTRIES>
                <ENTRY eventid="29" entrytime="00:01:20.82" heatid="29001" lane="4" />
                <ENTRY eventid="47" entrytime="00:01:20.29" heatid="47008" lane="2" />
                <ENTRY eventid="31" entrytime="00:01:11.91" heatid="31013" lane="1" />
                <ENTRY eventid="53" entrytime="00:02:54.37" heatid="53002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1506" eventid="29" swimtime="00:01:16.77" lane="4" heatid="29001" points="348">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1507" eventid="47" swimtime="00:01:16.95" lane="2" heatid="47008" points="362">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1508" eventid="31" swimtime="00:01:08.36" lane="1" heatid="31013" points="397">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1509" eventid="53" swimtime="00:02:52.43" lane="4" heatid="53002" points="352">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:18.52" />
                    <SPLIT distance="150" swimtime="00:02:10.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="338" birthdate="2015-01-01" gender="F" lastname="Treml" firstname="Lena" license="466283" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:47.87" heatid="3011" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:42.74" heatid="7013" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:44.81" heatid="9005" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:52.85" heatid="13003" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:41.70" heatid="15008" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:36.82" heatid="19010" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1510" eventid="3" swimtime="00:00:47.71" lane="4" heatid="3011" points="148" />
                <RESULT resultid="1511" eventid="7" swimtime="00:00:40.49" lane="4" heatid="7013" points="181" />
                <RESULT resultid="1512" eventid="9" swimtime="00:01:42.60" lane="2" heatid="9005" points="167">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1513" eventid="13" swimtime="00:00:50.65" lane="1" heatid="13003" points="111" />
                <RESULT resultid="1514" eventid="15" swimtime="00:01:42.44" lane="2" heatid="15008" points="153">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1515" eventid="19" swimtime="00:01:35.51" lane="1" heatid="19010" points="145">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="339" birthdate="2016-01-01" gender="F" lastname="Treml" firstname="Victoria" license="494868" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:53.78" heatid="3007" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:54.42" heatid="7004" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:55.00" heatid="9003" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:55.00" heatid="15005" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:45.00" heatid="19006" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1516" eventid="3" swimtime="00:00:53.11" lane="4" heatid="3007" points="107" />
                <RESULT resultid="1517" eventid="7" swimtime="00:00:55.77" lane="2" heatid="7004" points="69" />
                <RESULT resultid="1518" eventid="9" swimtime="00:02:07.93" lane="3" heatid="9003" points="86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1519" eventid="15" swimtime="00:01:59.59" lane="1" heatid="15005" points="96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1520" eventid="19" status="DSQ" swimtime="00:02:05.07" lane="3" heatid="19006" comment="Die Sportlerin startete vor dem Startsignal">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="340" birthdate="2004-01-01" gender="M" lastname="Walther" firstname="Theo" license="314090" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:26.06" heatid="44011" lane="3" />
                <ENTRY eventid="48" entrytime="00:01:03.40" heatid="48006" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:28.88" heatid="26006" lane="1" />
                <ENTRY eventid="32" entrytime="00:00:57.58" heatid="32009" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1521" eventid="44" swimtime="00:00:26.49" lane="3" heatid="44011" points="440" />
                <RESULT resultid="1522" eventid="48" swimtime="00:01:05.76" lane="3" heatid="48006" points="396">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1523" eventid="26" swimtime="00:00:29.61" lane="1" heatid="26006" points="416" />
                <RESULT resultid="1524" eventid="32" swimtime="00:00:58.03" lane="3" heatid="32009" points="461">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="341" birthdate="2015-01-01" gender="M" lastname="Weber" firstname="Fabien" license="466274">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:51.58" heatid="4004" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:41.41" heatid="8009" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:50.00" heatid="10002" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:50.00" heatid="16003" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:39.07" heatid="20005" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1525" eventid="4" swimtime="00:00:49.69" lane="3" heatid="4004" points="88" />
                <RESULT resultid="1526" eventid="8" swimtime="00:00:41.73" lane="1" heatid="8009" points="112" />
                <RESULT resultid="1527" eventid="10" swimtime="00:01:58.37" lane="3" heatid="10002" points="72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1528" eventid="16" swimtime="00:01:52.18" lane="4" heatid="16003" points="79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1529" eventid="20" swimtime="00:01:40.93" lane="1" heatid="20005" points="87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="342" birthdate="2017-01-01" gender="F" lastname="Zaiaieva" firstname="Dariia" license="496416" nation="UKR">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:02:05.07" heatid="5011" lane="1" />
                <ENTRY eventid="9" entrytime="00:02:00.00" heatid="9003" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:58.12" heatid="15005" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:59.62" heatid="17005" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:55.00" heatid="19004" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1530" eventid="5" swimtime="00:02:03.19" lane="1" heatid="5011" points="129">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1531" eventid="9" swimtime="00:02:04.53" lane="1" heatid="9003" points="93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1532" eventid="15" swimtime="00:01:57.08" lane="4" heatid="15005" points="103">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1533" eventid="17" swimtime="00:00:59.80" lane="3" heatid="17005" points="106" />
                <RESULT resultid="1534" eventid="19" swimtime="00:02:01.37" lane="4" heatid="19004" points="70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="343" birthdate="2013-01-01" gender="F" lastname="Zaiaieva" firstname="Vlada" license="468008" nation="UKR">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:33.43" heatid="1005" lane="1" />
                <ENTRY eventid="3" entrytime="00:00:35.85" heatid="3023" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:33.20" heatid="7030" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:25.21" heatid="9018" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:34.63" heatid="13016" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:19.32" heatid="15019" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1535" eventid="1" swimtime="00:01:27.98" lane="1" heatid="1005" points="231">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1536" eventid="3" swimtime="00:00:36.56" lane="3" heatid="3023" points="329" />
                <RESULT resultid="1537" eventid="7" swimtime="00:00:31.51" lane="3" heatid="7030" points="385" />
                <RESULT resultid="1538" eventid="9" swimtime="00:01:20.89" lane="4" heatid="9018" points="340">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1539" eventid="13" swimtime="00:00:34.45" lane="3" heatid="13016" points="354" />
                <RESULT resultid="1540" eventid="15" swimtime="00:01:22.62" lane="3" heatid="15019" points="293">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="344" birthdate="2014-01-01" gender="M" lastname="Zänsler" firstname="Elias" license="461989" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:39.52" heatid="2002" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:37.82" heatid="8012" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:35.00" heatid="10004" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:44.50" heatid="14005" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:24.92" heatid="20010" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1541" eventid="2" swimtime="00:01:36.43" lane="4" heatid="2002" points="121">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1542" eventid="8" swimtime="00:00:36.01" lane="1" heatid="8012" points="175" />
                <RESULT resultid="1543" eventid="10" swimtime="00:01:35.25" lane="3" heatid="10004" points="138">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1544" eventid="14" swimtime="00:00:44.24" lane="4" heatid="14005" points="118" />
                <RESULT resultid="1545" eventid="20" swimtime="00:01:22.99" lane="1" heatid="20010" points="157">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="345" birthdate="2014-01-01" gender="F" lastname="Zhokheieva" firstname="Mira" license="512067">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:48.01" heatid="3010" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:40.79" heatid="7015" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:45.00" heatid="13007" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:40.00" heatid="15009" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:25.00" heatid="19015" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1546" eventid="3" swimtime="00:00:47.48" lane="2" heatid="3010" points="150" />
                <RESULT resultid="1547" eventid="7" swimtime="00:00:40.71" lane="1" heatid="7015" points="178" />
                <RESULT resultid="1548" eventid="13" swimtime="00:00:44.82" lane="2" heatid="13007" points="160" />
                <RESULT resultid="1549" eventid="15" swimtime="00:01:52.03" lane="2" heatid="15009" points="117">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1550" eventid="19" swimtime="00:01:32.31" lane="3" heatid="19015" points="161">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="346" birthdate="2017-01-01" gender="F" lastname="Zhokheieva" firstname="Yuna" license="496417" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:50.32" heatid="3019" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:44.00" heatid="7026" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:50.57" heatid="9014" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:50.34" heatid="15015" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:43.55" heatid="19021" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1551" eventid="3" swimtime="00:00:48.06" lane="1" heatid="3019" points="145" />
                <RESULT resultid="1552" eventid="7" swimtime="00:00:44.50" lane="1" heatid="7026" points="136" />
                <RESULT resultid="1553" eventid="9" swimtime="00:01:49.27" lane="4" heatid="9014" points="138">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1554" eventid="15" swimtime="00:01:48.68" lane="2" heatid="15015" points="128">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1555" eventid="19" swimtime="00:01:40.42" lane="4" heatid="19021" points="125">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:41.82" lane="3" heatid="40003" />
                <ENTRY eventid="72" entrytime="00:01:51.03" lane="3" heatid="72003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1283" eventid="40" swimtime="00:01:36.56" lane="3" heatid="40003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.27" />
                    <SPLIT distance="100" swimtime="00:00:49.57" />
                    <SPLIT distance="150" swimtime="00:01:13.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="308" number="1" />
                    <RELAYPOSITION athleteid="331" number="2" />
                    <RELAYPOSITION athleteid="312" number="3" />
                    <RELAYPOSITION athleteid="328" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1284" eventid="72" swimtime="00:01:48.07" lane="3" heatid="72003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                    <SPLIT distance="100" swimtime="00:00:57.45" />
                    <SPLIT distance="150" swimtime="00:01:24.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="312" number="1" />
                    <RELAYPOSITION athleteid="331" number="2" />
                    <RELAYPOSITION athleteid="321" number="3" />
                    <RELAYPOSITION athleteid="328" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:02:04.55" lane="2" heatid="39001" />
                <ENTRY eventid="71" entrytime="00:02:12.06" lane="2" heatid="71002" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1285" eventid="39" swimtime="00:01:59.80" lane="2" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:00:58.75" />
                    <SPLIT distance="150" swimtime="00:01:29.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="310" number="1" />
                    <RELAYPOSITION athleteid="315" number="2" />
                    <RELAYPOSITION athleteid="337" number="3" />
                    <RELAYPOSITION athleteid="327" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1286" eventid="71" swimtime="00:02:10.01" lane="2" heatid="71002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="100" swimtime="00:01:07.25" />
                    <SPLIT distance="150" swimtime="00:01:39.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="315" number="1" />
                    <RELAYPOSITION athleteid="332" number="2" />
                    <RELAYPOSITION athleteid="311" number="3" />
                    <RELAYPOSITION athleteid="337" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:10.00" lane="2" heatid="11002" />
                <ENTRY eventid="23" entrytime="00:02:17.00" lane="2" heatid="23003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1287" eventid="11" swimtime="00:02:02.46" lane="2" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:02.29" />
                    <SPLIT distance="150" swimtime="00:01:30.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="343" number="1" />
                    <RELAYPOSITION athleteid="318" number="2" />
                    <RELAYPOSITION athleteid="332" number="3" />
                    <RELAYPOSITION athleteid="325" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1288" eventid="23" swimtime="00:02:15.60" lane="2" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:44.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="343" number="1" />
                    <RELAYPOSITION athleteid="318" number="2" />
                    <RELAYPOSITION athleteid="332" number="3" />
                    <RELAYPOSITION athleteid="325" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TJ Slávie Chomutov, z.s." nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="203" birthdate="2017-01-01" gender="F" lastname="BABKOVÁ" firstname="Katerina" license="63466969">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:58.51" heatid="3004" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:56.25" heatid="7003" lane="3" />
                <ENTRY eventid="17" entrytime="00:01:01.85" heatid="17004" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:53.90" heatid="19004" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="863" eventid="3" swimtime="00:00:57.07" lane="3" heatid="3004" points="86" />
                <RESULT resultid="864" eventid="7" swimtime="00:00:51.92" lane="3" heatid="7003" points="86" />
                <RESULT resultid="865" eventid="17" swimtime="00:00:59.41" lane="2" heatid="17004" points="108" />
                <RESULT resultid="866" eventid="19" swimtime="00:01:56.30" lane="1" heatid="19004" points="80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="204" birthdate="2016-01-01" gender="F" lastname="BELINGEROVÁ" firstname="Nikol" license="63455729">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.46" heatid="3020" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:36.17" heatid="7027" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:41.70" heatid="13013" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:20.88" heatid="19022" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="867" eventid="3" swimtime="00:00:41.70" lane="3" heatid="3020" points="222" />
                <RESULT resultid="868" eventid="7" swimtime="00:00:35.48" lane="1" heatid="7027" points="269" />
                <RESULT resultid="869" eventid="13" swimtime="00:00:39.66" lane="2" heatid="13013" points="232" />
                <RESULT resultid="870" eventid="19" swimtime="00:01:17.02" lane="2" heatid="19022" points="277">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="205" birthdate="2015-01-01" gender="F" lastname="BOROVICKOVÁ" firstname="Tereza" license="63471108">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:58.08" heatid="3005" lane="4" />
                <ENTRY eventid="5" entrytime="00:02:11.81" heatid="5003" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:46.49" heatid="7010" lane="4" />
                <ENTRY eventid="15" entrytime="00:02:01.94" heatid="15004" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:42.80" heatid="19008" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="871" eventid="3" swimtime="00:00:54.34" lane="4" heatid="3005" points="100" />
                <RESULT resultid="872" eventid="5" swimtime="00:02:10.67" lane="4" heatid="5003" points="108">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="873" eventid="7" swimtime="00:00:46.34" lane="4" heatid="7010" points="121" />
                <RESULT resultid="874" eventid="15" swimtime="00:01:58.69" lane="1" heatid="15004" points="98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="875" eventid="19" swimtime="00:01:41.31" lane="3" heatid="19008" points="122">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="206" birthdate="2017-01-01" gender="F" lastname="CERNEROVÁ" firstname="Hermína" license="63465407">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:52.41" heatid="3008" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:46.64" heatid="7026" lane="4" />
                <ENTRY eventid="17" entrytime="00:01:01.75" heatid="17005" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:41.28" heatid="19021" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="876" eventid="3" swimtime="00:00:48.30" lane="3" heatid="3008" points="142" />
                <RESULT resultid="877" eventid="7" swimtime="00:00:43.40" lane="4" heatid="7026" points="147" />
                <RESULT resultid="878" eventid="17" swimtime="00:01:00.68" lane="4" heatid="17005" points="102" />
                <RESULT resultid="879" eventid="19" swimtime="00:01:38.92" lane="1" heatid="19021" points="131">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="207" birthdate="2016-01-01" gender="F" lastname="CÍZKOVÁ" firstname="Adéla Ela" license="63471282">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:59.67" heatid="3003" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:59.38" heatid="7002" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:54.32" heatid="15005" lane="3" />
                <ENTRY eventid="17" entrytime="00:01:10.55" heatid="17003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="880" eventid="3" swimtime="00:01:04.14" lane="1" heatid="3003" points="61" />
                <RESULT resultid="881" eventid="7" swimtime="00:01:05.86" lane="1" heatid="7002" points="42" />
                <RESULT resultid="882" eventid="15" status="DSQ" swimtime="00:02:23.79" lane="3" heatid="15005" comment="Bei der zweiten Wende wurde die Wand nicht berührt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="883" eventid="17" status="DSQ" swimtime="00:01:02.44" lane="4" heatid="17003" comment="Die Sportlerin startete vor dem Startsignal" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="208" birthdate="2016-01-01" gender="F" lastname="CÍZKOVÁ" firstname="Anna Marie" license="63471283">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:54.47" heatid="3006" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:54.44" heatid="7004" lane="3" />
                <ENTRY eventid="17" entrytime="00:01:17.27" heatid="17002" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:44.49" heatid="19007" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="884" eventid="3" swimtime="00:00:53.20" lane="1" heatid="3006" points="106" />
                <RESULT resultid="885" eventid="7" swimtime="00:00:59.80" lane="3" heatid="7004" points="56" />
                <RESULT resultid="886" eventid="17" swimtime="00:01:08.66" lane="3" heatid="17002" points="70" />
                <RESULT resultid="887" eventid="19" swimtime="00:01:59.38" lane="1" heatid="19007" points="74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="209" birthdate="2014-01-01" gender="F" lastname="CÍZKOVÁ" firstname="Nela Eva" license="63458985">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:43.87" heatid="3015" lane="2" />
                <ENTRY eventid="5" entrytime="00:01:44.19" heatid="5008" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:37.17" heatid="7019" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:36.43" heatid="15010" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:48.87" heatid="17012" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:29.22" heatid="19014" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="888" eventid="3" swimtime="00:00:43.67" lane="2" heatid="3015" points="193" />
                <RESULT resultid="889" eventid="5" swimtime="00:01:47.40" lane="3" heatid="5008" points="195">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="890" eventid="7" swimtime="00:00:39.14" lane="3" heatid="7019" points="201" />
                <RESULT resultid="891" eventid="15" swimtime="00:01:37.09" lane="2" heatid="15010" points="180">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="892" eventid="17" swimtime="00:00:49.76" lane="4" heatid="17012" points="185" />
                <RESULT resultid="893" eventid="19" swimtime="00:01:33.62" lane="4" heatid="19014" points="154">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210" birthdate="2017-01-01" gender="F" lastname="CREPOVÁ" firstname="Karolína" license="63455732">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:44.85" heatid="3019" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:42.28" heatid="7026" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:59.44" heatid="17005" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:33.55" heatid="19021" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="894" eventid="3" swimtime="00:00:44.50" lane="2" heatid="3019" points="182" />
                <RESULT resultid="895" eventid="7" swimtime="00:00:40.71" lane="2" heatid="7026" points="178" />
                <RESULT resultid="896" eventid="17" swimtime="00:00:59.95" lane="2" heatid="17005" points="105" />
                <RESULT resultid="897" eventid="19" swimtime="00:01:32.69" lane="2" heatid="19021" points="159">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="211" birthdate="2016-01-01" gender="F" lastname="DOSTÁLOVÁ" firstname="Karla" license="63465386">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:59.06" heatid="3004" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:58.79" heatid="7002" lane="3" />
                <ENTRY eventid="17" entrytime="00:01:19.02" heatid="17002" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:43.83" heatid="19007" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="898" eventid="3" swimtime="00:01:05.78" lane="1" heatid="3004" points="56" />
                <RESULT resultid="899" eventid="7" swimtime="00:00:57.69" lane="3" heatid="7002" points="62" />
                <RESULT resultid="900" eventid="17" status="DSQ" swimtime="00:01:16.03" lane="1" heatid="17002" comment="Beim Zielanschlag hat die Sportlerin nicht mit beiden Händen gleichzeitig angeschlagen." />
                <RESULT resultid="901" eventid="19" swimtime="00:02:01.81" lane="2" heatid="19007" points="70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212" birthdate="2015-01-01" gender="M" lastname="FÁRA" firstname="Filip" license="63463229">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:46.31" heatid="4013" lane="3" />
                <ENTRY eventid="6" entrytime="00:02:05.43" heatid="6001" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:42.73" heatid="8008" lane="4" />
                <ENTRY eventid="16" entrytime="00:01:37.29" heatid="16008" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:39.06" heatid="20005" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="902" eventid="4" status="WDR" swimtime="00:00:00.00" lane="3" heatid="4013" />
                <RESULT resultid="903" eventid="6" status="WDR" swimtime="00:00:00.00" lane="2" heatid="6001" />
                <RESULT resultid="904" eventid="8" status="WDR" swimtime="00:00:00.00" lane="4" heatid="8008" />
                <RESULT resultid="905" eventid="16" status="WDR" swimtime="00:00:00.00" lane="3" heatid="16008" />
                <RESULT resultid="906" eventid="20" status="WDR" swimtime="00:00:00.00" lane="3" heatid="20005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213" birthdate="2014-01-01" gender="F" lastname="FEDERSELOVÁ" firstname="Ema" license="63445513">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:28.51" heatid="1004" lane="4" />
                <ENTRY eventid="5" entrytime="00:01:35.77" heatid="5010" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:26.01" heatid="9017" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:36.37" heatid="13015" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:22.03" heatid="15014" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:44.06" heatid="17019" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="907" eventid="1" swimtime="00:01:28.21" lane="4" heatid="1004" points="230">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="908" eventid="5" swimtime="00:01:38.16" lane="3" heatid="5010" points="256">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="909" eventid="9" swimtime="00:01:23.08" lane="4" heatid="9017" points="314">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="910" eventid="13" swimtime="00:00:36.29" lane="4" heatid="13015" points="303" />
                <RESULT resultid="911" eventid="15" swimtime="00:01:22.42" lane="2" heatid="15014" points="295">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="912" eventid="17" swimtime="00:00:43.91" lane="1" heatid="17019" points="269" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214" birthdate="2017-01-01" gender="F" lastname="FRICOVÁ" firstname="Barbora" license="63474210">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:02:06.39" heatid="5011" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:48.44" heatid="9014" lane="2" />
                <ENTRY eventid="13" entrytime="00:00:57.86" heatid="13012" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:55.80" heatid="17016" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="913" eventid="5" swimtime="00:01:58.25" lane="4" heatid="5011" points="146">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="914" eventid="9" swimtime="00:01:47.91" lane="2" heatid="9014" points="143">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="915" eventid="13" swimtime="00:00:56.23" lane="4" heatid="13012" points="81" />
                <RESULT resultid="916" eventid="17" swimtime="00:00:54.75" lane="1" heatid="17016" points="139" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="215" birthdate="2015-01-01" gender="M" lastname="GREGOR" firstname="Petr" license="63467320">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:51.94" heatid="4004" lane="4" />
                <ENTRY eventid="6" entrytime="00:01:51.54" heatid="6003" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:50.11" heatid="8004" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:53.38" heatid="18005" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:39.84" heatid="20004" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="917" eventid="4" status="WDR" swimtime="00:00:00.00" lane="4" heatid="4004" />
                <RESULT resultid="918" eventid="6" status="WDR" swimtime="00:00:00.00" lane="2" heatid="6003" />
                <RESULT resultid="919" eventid="8" status="WDR" swimtime="00:00:00.00" lane="4" heatid="8004" />
                <RESULT resultid="920" eventid="18" status="WDR" swimtime="00:00:00.00" lane="2" heatid="18005" />
                <RESULT resultid="921" eventid="20" status="WDR" swimtime="00:00:00.00" lane="2" heatid="20004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="216" birthdate="2017-01-01" gender="F" lastname="GREGOROVÁ" firstname="Barbara" license="63471154">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:53.02" heatid="3008" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:58.26" heatid="7002" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:58.92" heatid="15004" lane="2" />
                <ENTRY eventid="17" entrytime="00:01:20.28" heatid="17002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="922" eventid="3" swimtime="00:00:55.66" lane="4" heatid="3008" points="93" />
                <RESULT resultid="923" eventid="7" swimtime="00:00:54.48" lane="2" heatid="7002" points="74" />
                <RESULT resultid="924" eventid="15" status="DSQ" swimtime="00:02:01.74" lane="2" heatid="15004" comment="Die Sportlerin hat bei der zweiten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="925" eventid="17" status="DSQ" swimtime="00:01:09.96" lane="4" heatid="17002" comment="Beim Zielanschlag hat die Sportlerin nicht mit beiden Händen gleichzeitig angeschlagen." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="217" birthdate="2016-01-01" gender="M" lastname="HÁJEK" firstname="Josef" license="63460166">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:53.76" heatid="4003" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:42.44" heatid="8008" lane="1" />
                <ENTRY eventid="14" entrytime="00:01:00.59" heatid="14001" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:36.69" heatid="20006" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="926" eventid="4" swimtime="00:00:51.70" lane="1" heatid="4003" points="78" />
                <RESULT resultid="927" eventid="8" swimtime="00:00:42.21" lane="1" heatid="8008" points="108" />
                <RESULT resultid="928" eventid="14" swimtime="00:01:02.33" lane="2" heatid="14001" points="42" />
                <RESULT resultid="929" eventid="20" swimtime="00:01:37.43" lane="3" heatid="20006" points="97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="218" birthdate="2017-01-01" gender="F" lastname="HOLKOVÁ" firstname="Emma" license="63465359">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:54.73" heatid="3006" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:50.67" heatid="7006" lane="1" />
                <ENTRY eventid="17" entrytime="00:01:11.20" heatid="17002" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:52.16" heatid="19004" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="930" eventid="3" status="WDR" swimtime="00:00:00.00" lane="4" heatid="3006" />
                <RESULT resultid="931" eventid="7" status="WDR" swimtime="00:00:00.00" lane="1" heatid="7006" />
                <RESULT resultid="932" eventid="17" status="WDR" swimtime="00:00:00.00" lane="2" heatid="17002" />
                <RESULT resultid="933" eventid="19" status="WDR" swimtime="00:00:00.00" lane="3" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="219" birthdate="2014-01-01" gender="M" lastname="HOLÝ" firstname="Mikulás" license="63473213">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:39.18" heatid="4014" lane="4" />
                <ENTRY eventid="6" entrytime="00:01:46.98" heatid="6004" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:34.87" heatid="8015" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:45.94" heatid="14004" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:23.32" heatid="16009" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:16.24" heatid="20013" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="934" eventid="4" swimtime="00:00:36.82" lane="4" heatid="4014" points="216" />
                <RESULT resultid="935" eventid="6" swimtime="00:01:45.67" lane="2" heatid="6004" points="143">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="936" eventid="8" swimtime="00:00:33.53" lane="1" heatid="8015" points="217" />
                <RESULT resultid="937" eventid="14" swimtime="00:00:44.47" lane="2" heatid="14004" points="116" />
                <RESULT resultid="938" eventid="16" swimtime="00:01:22.10" lane="1" heatid="16009" points="203">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="939" eventid="20" swimtime="00:01:16.76" lane="2" heatid="20013" points="199">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="220" birthdate="2010-01-01" gender="M" lastname="JECMEN" firstname="Lukás" license="60117000">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:34.65" heatid="28005" lane="2" />
                <ENTRY eventid="38" entrytime="00:02:42.22" heatid="38005" lane="1" />
                <ENTRY eventid="46" entrytime="00:01:15.02" heatid="46003" lane="1" />
                <ENTRY eventid="54" entrytime="00:02:29.74" heatid="54003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="940" eventid="28" swimtime="00:00:34.44" lane="2" heatid="28005" points="380" />
                <RESULT resultid="941" eventid="38" swimtime="00:02:43.69" lane="1" heatid="38005" points="395">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:02:00.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="942" eventid="46" swimtime="00:01:15.58" lane="1" heatid="46003" points="391">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="943" eventid="54" swimtime="00:02:30.39" lane="4" heatid="54003" points="387">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                    <SPLIT distance="150" swimtime="00:01:54.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="221" birthdate="2010-01-01" gender="M" lastname="JECMEN" firstname="Petr" license="60118000">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:33.13" heatid="28007" lane="1" />
                <ENTRY eventid="38" entrytime="00:02:35.55" heatid="38006" lane="1" />
                <ENTRY eventid="46" entrytime="00:01:10.80" heatid="46005" lane="1" />
                <ENTRY eventid="54" entrytime="00:02:27.13" heatid="54003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="944" eventid="28" swimtime="00:00:32.78" lane="1" heatid="28007" points="440" />
                <RESULT resultid="945" eventid="38" swimtime="00:02:30.43" lane="1" heatid="38006" points="509">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="150" swimtime="00:01:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="946" eventid="46" swimtime="00:01:10.72" lane="1" heatid="46005" points="477">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="947" eventid="54" swimtime="00:02:27.10" lane="3" heatid="54003" points="413">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:13.69" />
                    <SPLIT distance="150" swimtime="00:01:52.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="222" birthdate="2007-01-01" gender="M" lastname="JEZBERA" firstname="Jakub" license="35718000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:26.79" heatid="44011" lane="4" />
                <ENTRY eventid="48" entrytime="00:00:59.47" heatid="48005" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:28.01" heatid="26009" lane="2" />
                <ENTRY eventid="36" entrytime="00:02:08.00" heatid="36003" lane="3" />
                <ENTRY eventid="54" entrytime="00:02:18.00" heatid="54005" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="948" eventid="44" swimtime="00:00:26.37" lane="4" heatid="44011" points="446" />
                <RESULT resultid="949" eventid="48" swimtime="00:00:59.46" lane="2" heatid="48005" points="537">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="950" eventid="26" swimtime="00:00:28.17" lane="2" heatid="26009" points="483" />
                <RESULT resultid="951" eventid="36" swimtime="00:02:09.87" lane="3" heatid="36003" points="538">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:03.00" />
                    <SPLIT distance="150" swimtime="00:01:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="952" eventid="54" swimtime="00:02:19.17" lane="1" heatid="54005" points="488">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                    <SPLIT distance="100" swimtime="00:01:06.13" />
                    <SPLIT distance="150" swimtime="00:01:47.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="223" birthdate="2015-01-01" gender="F" lastname="JURKOVÁ" firstname="Emma" license="63455737">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:51.88" heatid="3000" lane="0" />
                <ENTRY eventid="5" entrytime="00:02:14.20" heatid="5000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:45.35" heatid="7000" lane="0" />
                <ENTRY eventid="15" entrytime="00:01:48.28" heatid="15000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:43.96" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="953" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="954" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="955" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="956" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="957" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="224" birthdate="2014-01-01" gender="M" lastname="KARHAN" firstname="Kristián" license="63464637">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:34.18" heatid="6010" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:33.01" heatid="8019" lane="4" />
                <ENTRY eventid="10" entrytime="00:01:22.57" heatid="10011" lane="4" />
                <ENTRY eventid="16" entrytime="00:01:24.51" heatid="16009" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:44.06" heatid="18013" lane="2" />
                <ENTRY eventid="22" entrytime="00:02:55.90" heatid="22004" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="958" eventid="6" swimtime="00:01:30.00" lane="2" heatid="6010" points="231">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="959" eventid="8" swimtime="00:00:32.18" lane="4" heatid="8019" points="245" />
                <RESULT resultid="960" eventid="10" swimtime="00:01:21.60" lane="4" heatid="10011" points="220">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="961" eventid="16" status="DSQ" swimtime="00:01:22.50" lane="4" heatid="16009" comment="Der Sportler hat während der Schwimmstrecke die Rückenlage verlassen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="962" eventid="18" swimtime="00:00:41.45" lane="2" heatid="18013" points="218" />
                <RESULT resultid="963" eventid="22" swimtime="00:02:50.18" lane="1" heatid="22004" points="267">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:22.55" />
                    <SPLIT distance="150" swimtime="00:02:13.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="225" birthdate="2015-01-01" gender="F" lastname="KARHANOVÁ" firstname="Klaudie" license="63458975">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:38.49" heatid="1003" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:35.52" heatid="7023" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:26.31" heatid="9016" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:43.45" heatid="13009" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:25.62" heatid="15017" lane="2" />
                <ENTRY eventid="21" entrytime="00:03:07.69" heatid="21004" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="964" eventid="1" swimtime="00:01:36.44" lane="1" heatid="1003" points="176">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="965" eventid="7" swimtime="00:00:36.38" lane="3" heatid="7023" points="250" />
                <RESULT resultid="966" eventid="9" swimtime="00:01:29.63" lane="3" heatid="9016" points="250">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="967" eventid="13" swimtime="00:00:42.27" lane="4" heatid="13009" points="191" />
                <RESULT resultid="968" eventid="15" swimtime="00:01:27.49" lane="2" heatid="15017" points="246">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="969" eventid="21" swimtime="00:03:11.90" lane="4" heatid="21004" points="256">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                    <SPLIT distance="100" swimtime="00:01:34.87" />
                    <SPLIT distance="150" swimtime="00:02:29.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="226" birthdate="2010-01-01" gender="M" lastname="KOROUS" firstname="Matyás" license="60126000">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:32.28" heatid="28009" lane="1" />
                <ENTRY eventid="38" entrytime="00:02:28.94" heatid="38006" lane="3" />
                <ENTRY eventid="46" entrytime="00:01:10.22" heatid="46005" lane="3" />
                <ENTRY eventid="54" entrytime="00:02:19.39" heatid="54005" lane="4" />
                <ENTRY eventid="61" entrytime="00:00:31.98" heatid="61001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="970" eventid="28" swimtime="00:00:31.98" lane="1" heatid="28009" points="474" />
                <RESULT resultid="971" eventid="38" swimtime="00:02:28.31" lane="3" heatid="38006" points="531">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:12.53" />
                    <SPLIT distance="150" swimtime="00:01:50.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="972" eventid="46" swimtime="00:01:09.82" lane="3" heatid="46005" points="496">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="973" eventid="54" swimtime="00:02:18.58" lane="4" heatid="54005" points="495">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                    <SPLIT distance="150" swimtime="00:01:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2324" eventid="61" swimtime="00:00:31.84" lane="3" heatid="61001" points="481" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="227" birthdate="2014-01-01" gender="F" lastname="KOSTOLNÁ" firstname="Alice" license="63456889">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:38.12" heatid="3022" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:31.99" heatid="7029" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:27.66" heatid="9013" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:41.06" heatid="13010" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:18.27" heatid="15018" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:13.32" heatid="19024" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="974" eventid="3" status="WDR" swimtime="00:00:00.00" lane="3" heatid="3022" />
                <RESULT resultid="975" eventid="7" status="WDR" swimtime="00:00:00.00" lane="3" heatid="7029" />
                <RESULT resultid="976" eventid="9" status="WDR" swimtime="00:00:00.00" lane="4" heatid="9013" />
                <RESULT resultid="977" eventid="13" status="WDR" swimtime="00:00:00.00" lane="3" heatid="13010" />
                <RESULT resultid="978" eventid="15" status="WDR" swimtime="00:00:00.00" lane="2" heatid="15018">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="979" eventid="19" status="WDR" swimtime="00:00:00.00" lane="1" heatid="19024" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="228" birthdate="2013-01-01" gender="F" lastname="KREJCOVÁ" firstname="Viktorie" license="63455989">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:47.65" heatid="3011" lane="1" />
                <ENTRY eventid="5" entrytime="00:01:45.69" heatid="5007" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:39.06" heatid="7017" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:48.16" heatid="13005" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:49.50" heatid="17011" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:29.69" heatid="19013" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="980" eventid="3" swimtime="00:00:44.56" lane="1" heatid="3011" points="181" />
                <RESULT resultid="981" eventid="5" swimtime="00:01:44.48" lane="1" heatid="5007" points="212">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="982" eventid="7" swimtime="00:00:38.34" lane="3" heatid="7017" points="213" />
                <RESULT resultid="983" eventid="13" swimtime="00:00:46.50" lane="2" heatid="13005" points="144" />
                <RESULT resultid="984" eventid="17" swimtime="00:00:47.51" lane="2" heatid="17011" points="212" />
                <RESULT resultid="985" eventid="19" swimtime="00:01:29.27" lane="2" heatid="19013" points="178">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="229" birthdate="2008-01-01" gender="M" lastname="KUBISTA" firstname="Jan" license="58597000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:22.89" heatid="44000" lane="0" />
                <ENTRY eventid="34" entrytime="00:00:57.54" heatid="34000" lane="0" />
                <ENTRY eventid="42" entrytime="00:00:26.76" heatid="42000" lane="0" />
                <ENTRY eventid="26" entrytime="00:00:25.40" heatid="26000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="986" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="987" eventid="34" status="WDR" swimtime="00:00:00.00" lane="0" heatid="34000" />
                <RESULT resultid="988" eventid="42" status="WDR" swimtime="00:00:00.00" lane="0" heatid="42000" />
                <RESULT resultid="989" eventid="26" status="WDR" swimtime="00:00:00.00" lane="0" heatid="26000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="230" birthdate="2014-01-01" gender="M" lastname="KUNDRÁT" firstname="Jan" license="63462533">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:35.35" heatid="6010" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:31.99" heatid="8023" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:24.22" heatid="10007" lane="1" />
                <ENTRY eventid="14" entrytime="00:00:36.10" heatid="14010" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:44.36" heatid="18013" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:10.91" heatid="20020" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="990" eventid="6" swimtime="00:01:34.57" lane="3" heatid="6010" points="199">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="991" eventid="8" swimtime="00:00:30.95" lane="3" heatid="8023" points="276" />
                <RESULT resultid="992" eventid="10" swimtime="00:01:23.86" lane="1" heatid="10007" points="202">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="993" eventid="14" swimtime="00:00:37.13" lane="4" heatid="14010" points="201" />
                <RESULT resultid="994" eventid="18" swimtime="00:00:43.14" lane="3" heatid="18013" points="193" />
                <RESULT resultid="995" eventid="20" swimtime="00:01:09.84" lane="1" heatid="20020" points="264">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="231" birthdate="2015-01-01" gender="M" lastname="LEDEN" firstname="Teodor" license="63455744">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:41.96" heatid="2003" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:39.51" heatid="8011" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:38.78" heatid="10003" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:43.80" heatid="14009" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:54.98" heatid="18004" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:27.20" heatid="20009" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="996" eventid="2" swimtime="00:01:37.29" lane="2" heatid="2003" points="118">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="997" eventid="8" swimtime="00:00:36.95" lane="3" heatid="8011" points="162" />
                <RESULT resultid="998" eventid="10" swimtime="00:01:34.81" lane="3" heatid="10003" points="140">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="999" eventid="14" swimtime="00:00:44.55" lane="1" heatid="14009" points="116" />
                <RESULT resultid="1000" eventid="18" swimtime="00:00:53.43" lane="3" heatid="18004" points="101" />
                <RESULT resultid="1001" eventid="20" swimtime="00:01:25.03" lane="2" heatid="20009" points="146">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="232" birthdate="2016-01-01" gender="F" lastname="LEDNOVÁ" firstname="Laura" license="63455745">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:52.81" heatid="3008" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:48.00" heatid="7008" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:54.32" heatid="17007" lane="2" />
                <ENTRY eventid="19" entrytime="00:02:06.80" heatid="19002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1002" eventid="3" swimtime="00:00:51.77" lane="1" heatid="3008" points="116" />
                <RESULT resultid="1003" eventid="7" status="DSQ" swimtime="00:00:48.27" lane="2" heatid="7008" comment="Die Sportlerin startete vor dem Startsignal" />
                <RESULT resultid="1004" eventid="17" swimtime="00:01:03.75" lane="2" heatid="17007" points="88" />
                <RESULT resultid="1005" eventid="19" swimtime="00:01:45.68" lane="3" heatid="19002" points="107">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="233" birthdate="2010-01-01" gender="M" lastname="LICKO" firstname="Pavel" license="63436499">
              <ENTRIES>
                <ENTRY eventid="30" entrytime="00:01:03.57" heatid="30004" lane="4" />
                <ENTRY eventid="48" entrytime="00:01:02.65" heatid="48004" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:28.64" heatid="26008" lane="2" />
                <ENTRY eventid="36" entrytime="00:02:17.47" heatid="36003" lane="1" />
                <ENTRY eventid="57" entrytime="00:00:28.96" heatid="57001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1006" eventid="30" swimtime="00:01:04.71" lane="4" heatid="30004" points="402">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1007" eventid="48" swimtime="00:01:03.81" lane="2" heatid="48004" points="434">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1008" eventid="26" swimtime="00:00:28.96" lane="2" heatid="26008" points="445" />
                <RESULT resultid="1009" eventid="36" swimtime="00:02:19.82" lane="1" heatid="36003" points="431">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:09.24" />
                    <SPLIT distance="150" swimtime="00:01:45.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2358" eventid="57" swimtime="00:00:28.68" lane="4" heatid="57001" points="458" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="234" birthdate="2014-01-01" gender="F" lastname="MARKOVÁ" firstname="Nella" license="63450119">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:46.63" heatid="3013" lane="4" />
                <ENTRY eventid="5" entrytime="00:01:52.13" heatid="5006" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:40.57" heatid="7015" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:47.18" heatid="15007" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:53.15" heatid="17008" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:30.02" heatid="19013" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1010" eventid="3" swimtime="00:00:46.67" lane="4" heatid="3013" points="158" />
                <RESULT resultid="1011" eventid="5" swimtime="00:01:49.75" lane="4" heatid="5006" points="183">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1012" eventid="7" swimtime="00:00:41.19" lane="2" heatid="7015" points="172" />
                <RESULT resultid="1013" eventid="15" swimtime="00:01:43.26" lane="3" heatid="15007" points="150">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1014" eventid="17" swimtime="00:00:51.59" lane="3" heatid="17008" points="166" />
                <RESULT resultid="1015" eventid="19" swimtime="00:01:31.55" lane="3" heatid="19013" points="165">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="235" birthdate="2015-01-01" gender="M" lastname="MASOPUST" firstname="Mikulás" license="63456485">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:49.87" heatid="4000" lane="0" />
                <ENTRY eventid="6" entrytime="00:01:45.29" heatid="6000" lane="0" />
                <ENTRY eventid="8" entrytime="00:00:44.98" heatid="8000" lane="0" />
                <ENTRY eventid="16" entrytime="00:01:42.30" heatid="16000" lane="0" />
                <ENTRY eventid="18" entrytime="00:00:49.03" heatid="18000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1016" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="1017" eventid="6" status="WDR" swimtime="00:00:00.00" lane="0" heatid="6000" />
                <RESULT resultid="1018" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="1019" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="1020" eventid="18" status="WDR" swimtime="00:00:00.00" lane="0" heatid="18000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="236" birthdate="2014-01-01" gender="F" lastname="MATYSOVÁ" firstname="Klaudie" license="63480483">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:53.35" heatid="3007" lane="1" />
                <ENTRY eventid="5" entrytime="00:02:04.32" heatid="5003" lane="1" />
                <ENTRY eventid="7" entrytime="00:00:47.61" heatid="7009" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:53.17" heatid="15006" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:46.96" heatid="19006" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1021" eventid="3" swimtime="00:00:51.93" lane="1" heatid="3007" points="114" />
                <RESULT resultid="1022" eventid="5" swimtime="00:02:02.23" lane="1" heatid="5003" points="132">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1023" eventid="7" swimtime="00:00:45.37" lane="1" heatid="7009" points="129" />
                <RESULT resultid="1024" eventid="15" swimtime="00:01:56.70" lane="4" heatid="15006" points="104">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1025" eventid="19" swimtime="00:01:45.06" lane="4" heatid="19006" points="109">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="237" birthdate="2014-01-01" gender="F" lastname="MEINLOVÁ" firstname="Tereza" license="63445512">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:27.85" heatid="1004" lane="1" />
                <ENTRY eventid="5" entrytime="00:01:34.05" heatid="5014" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:25.23" heatid="9017" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:43.57" heatid="17019" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:15.02" heatid="19020" lane="3" />
                <ENTRY eventid="21" entrytime="00:02:59.31" heatid="21004" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1026" eventid="1" swimtime="00:01:32.99" lane="1" heatid="1004" points="196">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1027" eventid="5" swimtime="00:01:35.30" lane="4" heatid="5014" points="280">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1028" eventid="9" swimtime="00:01:27.25" lane="1" heatid="9017" points="271">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1029" eventid="17" swimtime="00:00:43.79" lane="3" heatid="17019" points="271" />
                <RESULT resultid="1030" eventid="19" swimtime="00:01:22.10" lane="3" heatid="19020" points="229">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1031" eventid="21" swimtime="00:03:09.24" lane="3" heatid="21004" points="267">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="100" swimtime="00:01:32.17" />
                    <SPLIT distance="150" swimtime="00:02:25.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="238" birthdate="2010-01-01" gender="M" lastname="MIKS" firstname="Ondrej" license="54734000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:26.32" heatid="44011" lane="1" />
                <ENTRY eventid="30" entrytime="00:01:02.96" heatid="30004" lane="3" />
                <ENTRY eventid="52" entrytime="00:02:02.25" heatid="52006" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:28.10" heatid="42011" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1032" eventid="44" swimtime="00:00:26.48" lane="1" heatid="44011" points="441" />
                <RESULT resultid="1033" eventid="30" swimtime="00:01:02.98" lane="3" heatid="30004" points="436">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1034" eventid="52" swimtime="00:02:04.56" lane="1" heatid="52006" points="507">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="100" swimtime="00:01:01.07" />
                    <SPLIT distance="150" swimtime="00:01:33.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1035" eventid="42" swimtime="00:00:28.02" lane="1" heatid="42011" points="467" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="239" birthdate="2015-01-01" gender="F" lastname="MIKSOVÁ" firstname="Ludmila" license="63455733">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:51.11" heatid="3000" lane="0" />
                <ENTRY eventid="5" entrytime="00:02:10.68" heatid="5000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:46.06" heatid="7000" lane="0" />
                <ENTRY eventid="15" entrytime="00:01:49.53" heatid="15000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:45.16" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1036" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="1037" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="1038" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="1039" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="1040" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="240" birthdate="2007-01-01" gender="F" lastname="NEVOLOVÁ" firstname="Katerina" license="45348000">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:29.86" heatid="43013" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:09.66" heatid="47007" lane="2" />
                <ENTRY eventid="25" entrytime="00:00:33.13" heatid="25008" lane="2" />
                <ENTRY eventid="49" entrytime="00:02:43.64" heatid="49001" lane="1" />
                <ENTRY eventid="35" entrytime="00:02:30.05" heatid="35003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1041" eventid="43" swimtime="00:00:29.57" lane="3" heatid="43013" points="466" />
                <RESULT resultid="1042" eventid="47" swimtime="00:01:10.26" lane="2" heatid="47007" points="476">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1043" eventid="25" swimtime="00:00:32.70" lane="2" heatid="25008" points="460" />
                <RESULT resultid="1044" eventid="49" swimtime="00:02:38.33" lane="1" heatid="49001" points="431">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:14.74" />
                    <SPLIT distance="150" swimtime="00:01:56.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1045" eventid="35" swimtime="00:02:33.01" lane="3" heatid="35003" points="469">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:15.00" />
                    <SPLIT distance="150" swimtime="00:01:54.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="241" birthdate="2016-01-01" gender="M" lastname="NGUYEN DANG" firstname="Gia Hao" license="63458977">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:51.55" heatid="4004" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:43.32" heatid="8007" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:57.52" heatid="18003" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:38.36" heatid="20005" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1046" eventid="4" status="WDR" swimtime="00:00:00.00" lane="2" heatid="4004" />
                <RESULT resultid="1047" eventid="8" status="WDR" swimtime="00:00:00.00" lane="1" heatid="8007" />
                <RESULT resultid="1048" eventid="18" status="WDR" swimtime="00:00:00.00" lane="3" heatid="18003" />
                <RESULT resultid="1049" eventid="20" status="WDR" swimtime="00:00:00.00" lane="2" heatid="20005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="242" birthdate="2015-01-01" gender="F" lastname="NGUYEN" firstname="Ella" license="63455748">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:47.64" heatid="3011" lane="3" />
                <ENTRY eventid="5" entrytime="00:01:55.45" heatid="5005" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:38.97" heatid="7017" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:39.00" heatid="15010" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:53.36" heatid="17008" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:24.28" heatid="19015" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1050" eventid="3" swimtime="00:00:48.15" lane="3" heatid="3011" points="144" />
                <RESULT resultid="1051" eventid="5" swimtime="00:01:52.16" lane="4" heatid="5005" points="171">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1052" eventid="7" swimtime="00:00:38.12" lane="2" heatid="7017" points="217" />
                <RESULT resultid="1053" eventid="15" swimtime="00:01:41.76" lane="1" heatid="15010" points="156">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1054" eventid="17" swimtime="00:00:52.89" lane="1" heatid="17008" points="154" />
                <RESULT resultid="1055" eventid="19" swimtime="00:01:28.74" lane="2" heatid="19015" points="181">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="243" birthdate="2017-01-01" gender="M" lastname="PECHÁC" firstname="David" license="63458970">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:55.23" heatid="4011" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:52.80" heatid="8003" lane="1" />
                <ENTRY eventid="18" entrytime="00:01:20.15" heatid="18001" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:54.51" heatid="20003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1056" eventid="4" swimtime="00:00:56.87" lane="3" heatid="4011" points="58" />
                <RESULT resultid="1057" eventid="8" swimtime="00:00:53.21" lane="1" heatid="8003" points="54" />
                <RESULT resultid="1058" eventid="18" swimtime="00:01:18.28" lane="3" heatid="18001" points="32" />
                <RESULT resultid="1059" eventid="20" swimtime="00:02:01.94" lane="4" heatid="20003" points="49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="244" birthdate="2009-01-01" gender="M" lastname="PECHÁC" firstname="Denis" license="54739000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:29.32" heatid="44005" lane="3" />
                <ENTRY eventid="34" entrytime="00:01:14.80" heatid="34004" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:34.47" heatid="42003" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:34.20" heatid="26003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1060" eventid="44" swimtime="00:00:28.41" lane="3" heatid="44005" points="357" />
                <RESULT resultid="1061" eventid="34" swimtime="00:01:13.64" lane="3" heatid="34004" points="299">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1062" eventid="42" swimtime="00:00:34.29" lane="2" heatid="42003" points="255" />
                <RESULT resultid="1063" eventid="26" swimtime="00:00:33.23" lane="2" heatid="26003" points="294" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="245" birthdate="2014-01-01" gender="M" lastname="ROUC" firstname="Vlastimil" license="63467317">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:22.40" heatid="2004" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:32.18" heatid="8023" lane="1" />
                <ENTRY eventid="10" entrytime="00:01:24.16" heatid="10007" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:35.71" heatid="14010" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:11.37" heatid="20020" lane="4" />
                <ENTRY eventid="22" entrytime="00:02:58.60" heatid="22004" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1064" eventid="2" swimtime="00:01:18.75" lane="3" heatid="2004" points="223">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1065" eventid="8" swimtime="00:00:30.85" lane="1" heatid="8023" points="279" />
                <RESULT resultid="1066" eventid="10" swimtime="00:01:21.34" lane="3" heatid="10007" points="222">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1067" eventid="14" swimtime="00:00:34.47" lane="1" heatid="14010" points="251" />
                <RESULT resultid="1068" eventid="20" swimtime="00:01:07.73" lane="4" heatid="20020" points="290">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1069" eventid="22" swimtime="00:02:49.14" lane="4" heatid="22004" points="272">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:21.33" />
                    <SPLIT distance="150" swimtime="00:02:13.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="246" birthdate="2008-01-01" gender="M" lastname="ROUS" firstname="David" license="42028000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.95" heatid="44016" lane="4" />
                <ENTRY eventid="48" entrytime="00:01:00.80" heatid="48005" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:28.62" heatid="26009" lane="4" />
                <ENTRY eventid="32" entrytime="00:00:54.71" heatid="32012" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1070" eventid="44" status="WDR" swimtime="00:00:00.00" lane="4" heatid="44016" />
                <RESULT resultid="1071" eventid="48" status="WDR" swimtime="00:00:00.00" lane="3" heatid="48005" />
                <RESULT resultid="1072" eventid="26" status="WDR" swimtime="00:00:00.00" lane="4" heatid="26009" />
                <RESULT resultid="1073" eventid="32" status="WDR" swimtime="00:00:00.00" lane="4" heatid="32012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="247" birthdate="2015-01-01" gender="F" lastname="RUZKOVÁ" firstname="Ella" license="63447073">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:36.02" heatid="1003" lane="3" />
                <ENTRY eventid="3" entrytime="00:00:43.07" heatid="3016" lane="3" />
                <ENTRY eventid="9" entrytime="00:01:29.81" heatid="9016" lane="1" />
                <ENTRY eventid="13" entrytime="00:00:39.22" heatid="13014" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:17.59" heatid="19023" lane="3" />
                <ENTRY eventid="21" entrytime="00:03:12.70" heatid="21003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1074" eventid="1" swimtime="00:01:39.68" lane="3" heatid="1003" points="159">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1075" eventid="3" swimtime="00:00:44.35" lane="3" heatid="3016" points="184" />
                <RESULT resultid="1076" eventid="9" swimtime="00:01:29.50" lane="1" heatid="9016" points="251">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1077" eventid="13" swimtime="00:00:39.67" lane="2" heatid="13014" points="232" />
                <RESULT resultid="1078" eventid="19" swimtime="00:01:18.76" lane="3" heatid="19023" points="259">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1079" eventid="21" swimtime="00:03:22.77" lane="1" heatid="21003" points="217">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                    <SPLIT distance="100" swimtime="00:01:38.50" />
                    <SPLIT distance="150" swimtime="00:02:37.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="248" birthdate="2013-01-01" gender="M" lastname="RYBÁR" firstname="Matej" license="63481090">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:55.11" heatid="4002" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:44.75" heatid="8005" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:54.21" heatid="16002" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:48.78" heatid="20003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1080" eventid="4" swimtime="00:00:51.68" lane="2" heatid="4002" points="78" />
                <RESULT resultid="1081" eventid="8" swimtime="00:00:41.14" lane="2" heatid="8005" points="117" />
                <RESULT resultid="1082" eventid="16" swimtime="00:01:52.60" lane="2" heatid="16002" points="79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1083" eventid="20" swimtime="00:01:36.82" lane="3" heatid="20003" points="99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="249" birthdate="2017-01-01" gender="F" lastname="RYBÁROVÁ" firstname="Johanka" license="63471886">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:59.83" heatid="3003" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:56.74" heatid="7003" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:59.16" heatid="15004" lane="3" />
                <ENTRY eventid="17" entrytime="00:01:24.97" heatid="17001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1084" eventid="3" swimtime="00:00:58.75" lane="4" heatid="3003" points="79" />
                <RESULT resultid="1085" eventid="7" swimtime="00:00:59.26" lane="1" heatid="7003" points="57" />
                <RESULT resultid="1086" eventid="15" swimtime="00:02:17.92" lane="3" heatid="15004" points="63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1087" eventid="17" swimtime="00:01:14.89" lane="2" heatid="17001" points="54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="250" birthdate="2015-01-01" gender="F" lastname="SCHNITTEROVÁ" firstname="Adéla" license="63458976">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:41.63" heatid="5013" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:36.31" heatid="7021" lane="2" />
                <ENTRY eventid="9" entrytime="00:01:30.23" heatid="9012" lane="4" />
                <ENTRY eventid="13" entrytime="00:00:43.54" heatid="13008" lane="2" />
                <ENTRY eventid="15" entrytime="00:01:28.33" heatid="15017" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:21.95" heatid="19018" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1088" eventid="5" swimtime="00:01:40.69" lane="4" heatid="5013" points="237">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1089" eventid="7" swimtime="00:00:37.27" lane="2" heatid="7021" points="232" />
                <RESULT resultid="1090" eventid="9" swimtime="00:01:30.89" lane="4" heatid="9012" points="240">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1091" eventid="13" status="DNS" swimtime="00:00:00.00" lane="2" heatid="13008" />
                <RESULT resultid="1092" eventid="15" status="DNS" swimtime="00:00:00.00" lane="4" heatid="15017" />
                <RESULT resultid="1093" eventid="19" status="DNS" swimtime="00:00:00.00" lane="3" heatid="19018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="251" birthdate="2008-01-01" gender="M" lastname="SELINGR" firstname="Lukás" license="49585000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:23.80" heatid="44016" lane="2" />
                <ENTRY eventid="30" entrytime="00:00:55.05" heatid="30005" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:25.13" heatid="42012" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:28.48" heatid="26009" lane="1" />
                <ENTRY eventid="32" entrytime="00:00:52.49" heatid="32012" lane="2" />
                <ENTRY eventid="69" entrytime="00:00:25.15" heatid="69001" lane="4" />
                <ENTRY eventid="66" entrytime="00:00:25.54" heatid="66001" lane="1" />
                <ENTRY eventid="57" entrytime="00:00:28.18" heatid="57001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1094" eventid="44" swimtime="00:00:25.15" lane="2" heatid="44016" points="515" />
                <RESULT resultid="1095" eventid="30" swimtime="00:00:58.01" lane="2" heatid="30005" points="558">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1096" eventid="42" swimtime="00:00:25.54" lane="2" heatid="42012" points="617" />
                <RESULT resultid="1097" eventid="26" swimtime="00:00:28.18" lane="1" heatid="26009" points="482" />
                <RESULT resultid="1098" eventid="32" swimtime="00:00:54.21" lane="2" heatid="32012" points="565">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2356" eventid="57" swimtime="00:00:27.53" lane="3" heatid="57001" points="518" />
                <RESULT resultid="2345" eventid="66" swimtime="00:00:25.53" lane="1" heatid="66001" points="618" />
                <RESULT resultid="2310" eventid="69" swimtime="00:00:24.91" lane="4" heatid="69001" points="530" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="252" birthdate="2010-01-01" gender="F" lastname="SILNÁ" firstname="Barbora" license="56500000">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:35.67" heatid="27008" lane="3" />
                <ENTRY eventid="33" entrytime="00:01:10.02" heatid="33008" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:30.69" heatid="41010" lane="1" />
                <ENTRY eventid="45" entrytime="00:01:16.31" heatid="45006" lane="2" />
                <ENTRY eventid="59" entrytime="00:00:36.76" heatid="59001" lane="3" />
                <ENTRY eventid="63" entrytime="00:00:31.48" heatid="63001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1099" eventid="27" swimtime="00:00:36.76" lane="3" heatid="27008" points="459" />
                <RESULT resultid="1100" eventid="33" swimtime="00:01:11.28" lane="3" heatid="33008" points="498">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1101" eventid="41" swimtime="00:00:31.48" lane="1" heatid="41010" points="464" />
                <RESULT resultid="1102" eventid="45" swimtime="00:01:18.25" lane="2" heatid="45006" points="506">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2316" eventid="59" swimtime="00:00:35.57" lane="3" heatid="59001" points="507" />
                <RESULT resultid="2332" eventid="63" swimtime="00:00:31.22" lane="3" heatid="63001" points="476" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="253" birthdate="2014-01-01" gender="F" lastname="SLÁDECKOVÁ" firstname="Lea" license="63465404">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:23.67" heatid="1004" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:33.34" heatid="7029" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:24.96" heatid="9017" lane="3" />
                <ENTRY eventid="13" entrytime="00:00:35.50" heatid="13015" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:20.97" heatid="15018" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:11.97" heatid="19024" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1103" eventid="1" swimtime="00:01:24.33" lane="3" heatid="1004" points="263">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1104" eventid="7" swimtime="00:00:33.57" lane="4" heatid="7029" points="318" />
                <RESULT resultid="1105" eventid="9" swimtime="00:01:22.96" lane="3" heatid="9017" points="316">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1106" eventid="13" swimtime="00:00:36.35" lane="3" heatid="13015" points="301" />
                <RESULT resultid="1107" eventid="15" swimtime="00:01:21.28" lane="4" heatid="15018" points="307">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1108" eventid="19" swimtime="00:01:12.90" lane="3" heatid="19024" points="327">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="254" birthdate="2009-01-01" gender="F" lastname="STANKOVÁ" firstname="Katerina" license="49588000">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:29.55" heatid="43008" lane="2" />
                <ENTRY eventid="47" entrytime="00:01:07.16" heatid="47006" lane="2" />
                <ENTRY eventid="25" entrytime="00:00:31.57" heatid="25007" lane="1" />
                <ENTRY eventid="35" entrytime="00:02:29.16" heatid="35003" lane="2" />
                <ENTRY eventid="67" entrytime="00:00:29.28" heatid="67001" lane="4" />
                <ENTRY eventid="56" entrytime="00:00:31.95" heatid="56001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1109" eventid="43" swimtime="00:00:29.28" lane="2" heatid="43008" points="480" />
                <RESULT resultid="1110" eventid="47" swimtime="00:01:07.83" lane="2" heatid="47006" points="529">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1111" eventid="25" swimtime="00:00:31.95" lane="1" heatid="25007" points="493" />
                <RESULT resultid="1112" eventid="35" swimtime="00:02:25.65" lane="2" heatid="35003" points="544">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:11.45" />
                    <SPLIT distance="150" swimtime="00:01:48.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2353" eventid="56" swimtime="00:00:31.97" lane="1" heatid="56001" points="492" />
                <RESULT resultid="2302" eventid="67" swimtime="00:00:29.01" lane="4" heatid="67001" points="493" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="255" birthdate="2010-01-01" gender="M" lastname="STUDENT" firstname="Tobias" license="49783000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:25.07" heatid="44015" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:31.66" heatid="28009" lane="3" />
                <ENTRY eventid="34" entrytime="00:00:59.78" heatid="34007" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:27.16" heatid="42011" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:29.36" heatid="26008" lane="3" />
                <ENTRY eventid="69" entrytime="00:00:24.74" heatid="69001" lane="2" />
                <ENTRY eventid="61" entrytime="00:00:30.95" heatid="61001" lane="2" />
                <ENTRY eventid="65" entrytime="00:00:26.80" heatid="65001" lane="3" />
                <ENTRY eventid="57" entrytime="00:00:27.65" heatid="57001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1113" eventid="44" swimtime="00:00:24.74" lane="2" heatid="44015" points="541" />
                <RESULT resultid="1114" eventid="28" swimtime="00:00:30.95" lane="3" heatid="28009" points="523" />
                <RESULT resultid="1115" eventid="34" swimtime="00:00:59.59" lane="2" heatid="34007" points="565">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1116" eventid="42" swimtime="00:00:26.80" lane="3" heatid="42011" points="534" />
                <RESULT resultid="1117" eventid="26" swimtime="00:00:27.65" lane="3" heatid="26008" points="511" />
                <RESULT resultid="2355" eventid="57" swimtime="00:00:27.43" lane="2" heatid="57001" points="523" />
                <RESULT resultid="2323" eventid="61" swimtime="00:00:31.02" lane="2" heatid="61001" points="520" />
                <RESULT resultid="2340" eventid="65" swimtime="00:00:26.83" lane="3" heatid="65001" points="532" />
                <RESULT resultid="2307" eventid="69" swimtime="00:00:25.00" lane="2" heatid="69001" points="524" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="256" birthdate="2010-01-01" gender="M" lastname="STUDNICKA" firstname="Simon" license="54758000">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:29.68" heatid="28009" lane="2" />
                <ENTRY eventid="38" entrytime="00:02:16.34" heatid="38006" lane="2" />
                <ENTRY eventid="46" entrytime="00:01:03.05" heatid="46005" lane="2" />
                <ENTRY eventid="54" entrytime="00:02:06.26" heatid="54005" lane="2" />
                <ENTRY eventid="62" entrytime="00:00:29.48" heatid="62001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1118" eventid="28" swimtime="00:00:29.48" lane="2" heatid="28009" points="606" />
                <RESULT resultid="1119" eventid="38" swimtime="00:02:21.57" lane="2" heatid="38006" points="611">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:45.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1120" eventid="46" swimtime="00:01:03.87" lane="2" heatid="46005" points="648">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1121" eventid="54" swimtime="00:02:10.03" lane="2" heatid="54005" points="599">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="100" swimtime="00:01:02.68" />
                    <SPLIT distance="150" swimtime="00:01:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2328" eventid="62" swimtime="00:00:29.44" lane="3" heatid="62001" points="608" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="257" birthdate="2010-01-01" gender="F" lastname="SURKOVÁ" firstname="Barbora" license="63438636">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:26.51" heatid="43012" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:34.49" heatid="27008" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:07.91" heatid="33008" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:30.20" heatid="41010" lane="3" />
                <ENTRY eventid="31" entrytime="00:00:59.47" heatid="31011" lane="2" />
                <ENTRY eventid="68" entrytime="00:00:26.69" heatid="68001" lane="3" />
                <ENTRY eventid="60" entrytime="00:00:34.24" heatid="60001" lane="3" />
                <ENTRY eventid="64" entrytime="00:00:30.22" heatid="64001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1122" eventid="43" swimtime="00:00:26.69" lane="3" heatid="43012" points="634" />
                <RESULT resultid="1123" eventid="27" swimtime="00:00:34.24" lane="2" heatid="27008" points="568" />
                <RESULT resultid="1124" eventid="33" swimtime="00:01:09.39" lane="2" heatid="33008" points="540">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1125" eventid="41" swimtime="00:00:30.22" lane="3" heatid="41010" points="525" />
                <RESULT resultid="1126" eventid="31" swimtime="00:01:00.82" lane="2" heatid="31011" points="563">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2320" eventid="60" swimtime="00:00:33.58" lane="3" heatid="60001" points="603" />
                <RESULT resultid="2336" eventid="64" swimtime="00:00:30.15" lane="3" heatid="64001" points="528" />
                <RESULT resultid="2304" eventid="68" swimtime="00:00:26.37" lane="3" heatid="68001" points="657" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="258" birthdate="2010-01-01" gender="M" lastname="SÝKORA" firstname="Jakub" license="57945000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.64" heatid="44008" lane="4" />
                <ENTRY eventid="48" entrytime="00:01:04.81" heatid="48004" lane="3" />
                <ENTRY eventid="50" entrytime="00:02:18.74" heatid="50002" lane="3" />
                <ENTRY eventid="54" entrytime="00:02:19.64" heatid="54004" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1127" eventid="44" swimtime="00:00:27.29" lane="4" heatid="44008" points="403" />
                <RESULT resultid="1128" eventid="48" swimtime="00:01:04.18" lane="3" heatid="48004" points="427">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1129" eventid="50" swimtime="00:02:20.18" lane="3" heatid="50002" points="442">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:06.27" />
                    <SPLIT distance="150" swimtime="00:01:43.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1130" eventid="54" swimtime="00:02:19.30" lane="2" heatid="54004" points="487">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="100" swimtime="00:01:04.97" />
                    <SPLIT distance="150" swimtime="00:01:46.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="259" birthdate="2007-01-01" gender="F" lastname="VLASÁKOVÁ" firstname="Tereza" license="45354000">
              <ENTRIES>
                <ENTRY eventid="29" entrytime="00:01:05.20" heatid="29006" lane="2" />
                <ENTRY eventid="37" entrytime="00:02:47.10" heatid="37002" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:30.10" heatid="41011" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:16.50" heatid="45007" lane="3" />
                <ENTRY eventid="49" entrytime="00:02:26.50" heatid="49001" lane="2" />
                <ENTRY eventid="64" entrytime="00:00:30.30" heatid="64001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1131" eventid="29" swimtime="00:01:07.06" lane="2" heatid="29006" points="523">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1132" eventid="37" swimtime="00:02:46.97" lane="1" heatid="37002" points="523">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:20.13" />
                    <SPLIT distance="150" swimtime="00:02:03.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1133" eventid="41" swimtime="00:00:30.30" lane="2" heatid="41011" points="520" />
                <RESULT resultid="1134" eventid="45" swimtime="00:01:17.51" lane="3" heatid="45007" points="520">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1135" eventid="49" swimtime="00:02:33.95" lane="2" heatid="49001" points="468">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2337" eventid="64" swimtime="00:00:30.07" lane="1" heatid="64001" points="532" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="260" birthdate="2010-01-01" gender="M" lastname="VOKATÝ" firstname="Matej" license="60186000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:25.08" heatid="44015" lane="3" />
                <ENTRY eventid="52" entrytime="00:02:01.51" heatid="52006" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:28.63" heatid="42007" lane="1" />
                <ENTRY eventid="32" entrytime="00:00:55.39" heatid="32011" lane="2" />
                <ENTRY eventid="69" entrytime="00:00:24.95" heatid="69001" lane="1" />
                <ENTRY eventid="65" entrytime="00:00:27.90" heatid="65001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1136" eventid="44" swimtime="00:00:24.95" lane="3" heatid="44015" points="527" />
                <RESULT resultid="1137" eventid="52" swimtime="00:02:03.01" lane="3" heatid="52006" points="527">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="100" swimtime="00:00:58.84" />
                    <SPLIT distance="150" swimtime="00:01:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1138" eventid="42" swimtime="00:00:27.90" lane="1" heatid="42007" points="473" />
                <RESULT resultid="1139" eventid="32" swimtime="00:00:55.43" lane="2" heatid="32011" points="529">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2342" eventid="65" swimtime="00:00:27.69" lane="4" heatid="65001" points="484" />
                <RESULT resultid="2309" eventid="69" swimtime="00:00:24.97" lane="1" heatid="69001" points="526" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="261" birthdate="2014-01-01" gender="M" lastname="VURBS" firstname="Ondrej" license="63455754">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:27.51" heatid="2004" lane="4" />
                <ENTRY eventid="4" entrytime="00:00:40.72" heatid="4010" lane="3" />
                <ENTRY eventid="10" entrytime="00:01:28.00" heatid="10006" lane="3" />
                <ENTRY eventid="14" entrytime="00:00:38.23" heatid="14006" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:26.66" heatid="16005" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:15.42" heatid="20014" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1140" eventid="2" swimtime="00:01:28.96" lane="4" heatid="2004" points="154">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1141" eventid="4" swimtime="00:00:40.75" lane="3" heatid="4010" points="159" />
                <RESULT resultid="1142" eventid="10" swimtime="00:01:25.57" lane="3" heatid="10006" points="191">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1143" eventid="14" swimtime="00:00:36.75" lane="2" heatid="14006" points="207" />
                <RESULT resultid="1144" eventid="16" swimtime="00:01:27.63" lane="2" heatid="16005" points="167">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1145" eventid="20" swimtime="00:01:14.63" lane="1" heatid="20014" points="216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="262" birthdate="2013-01-01" gender="F" lastname="ZÁRECKÁ" firstname="Ella" license="63455833">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:58.79" heatid="3000" lane="0" />
                <ENTRY eventid="5" entrytime="00:02:19.55" heatid="5000" lane="0" />
                <ENTRY eventid="7" entrytime="00:00:48.17" heatid="7000" lane="0" />
                <ENTRY eventid="15" entrytime="00:02:07.95" heatid="15000" lane="0" />
                <ENTRY eventid="19" entrytime="00:01:51.05" heatid="19000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1146" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="1147" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="1148" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="1149" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="1150" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="263" birthdate="2015-01-01" gender="M" lastname="ZÁRECKÝ" firstname="Dan" license="63455832">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:53.57" heatid="4000" lane="0" />
                <ENTRY eventid="6" entrytime="00:02:05.79" heatid="6000" lane="0" />
                <ENTRY eventid="8" entrytime="00:00:47.88" heatid="8000" lane="0" />
                <ENTRY eventid="16" entrytime="00:01:54.12" heatid="16000" lane="0" />
                <ENTRY eventid="18" entrytime="00:00:55.11" heatid="18000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1151" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="1152" eventid="6" status="WDR" swimtime="00:00:00.00" lane="0" heatid="6000" />
                <RESULT resultid="1153" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="1154" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="1155" eventid="18" status="WDR" swimtime="00:00:00.00" lane="0" heatid="18000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="493" birthdate="2012-01-01" gender="F" lastname="Kvetová" firstname="Markéta" license="0">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:40.68" heatid="27006" lane="1" />
                <ENTRY eventid="29" entrytime="00:01:29.58" heatid="29002" lane="1" />
                <ENTRY eventid="37" entrytime="00:03:08.67" heatid="37001" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:28.10" heatid="45004" lane="2" />
                <ENTRY eventid="53" entrytime="00:02:55.06" heatid="53001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2274" eventid="27" swimtime="00:00:41.24" lane="1" heatid="27006" points="325" />
                <RESULT resultid="2275" eventid="29" swimtime="00:01:32.75" lane="1" heatid="29002" points="197">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2276" eventid="37" swimtime="00:03:09.49" lane="2" heatid="37001" points="358">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:32.20" />
                    <SPLIT distance="150" swimtime="00:02:22.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2277" eventid="45" swimtime="00:01:29.05" lane="2" heatid="45004" points="343">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2278" eventid="53" swimtime="00:02:54.57" lane="3" heatid="53001" points="340">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:14.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="494" birthdate="2012-01-01" gender="M" lastname="Masopust" firstname="Tomás" license="0" nation="CZE">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:01:17.38" heatid="10013" lane="2" />
                <ENTRY eventid="16" entrytime="00:01:20.11" heatid="16011" lane="2" />
                <ENTRY eventid="22" entrytime="00:02:46.50" heatid="22005" lane="1" />
                <ENTRY eventid="6" entrytime="00:01:25.84" heatid="6012" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:33.19" heatid="8018" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2279" eventid="6" swimtime="00:01:25.65" lane="1" heatid="6012" points="268">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2280" eventid="8" swimtime="00:00:33.03" lane="4" heatid="8018" points="227" />
                <RESULT resultid="2281" eventid="10" swimtime="00:01:18.10" lane="2" heatid="10013" points="251">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2282" eventid="16" swimtime="00:01:18.26" lane="2" heatid="16011" points="235">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2283" eventid="22" swimtime="00:02:48.07" lane="1" heatid="22005" points="277">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                    <SPLIT distance="100" swimtime="00:01:19.97" />
                    <SPLIT distance="150" swimtime="00:02:09.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="495" birthdate="2011-01-01" gender="M" lastname="Hrych" firstname="Jan" license="0">
              <ENTRIES>
                <ENTRY eventid="36" entrytime="00:02:29.35" heatid="36002" lane="3" />
                <ENTRY eventid="44" entrytime="00:00:29.38" heatid="44014" lane="1" />
                <ENTRY eventid="48" entrytime="00:01:08.96" heatid="48003" lane="2" />
                <ENTRY eventid="52" entrytime="00:02:19.68" heatid="52004" lane="3" />
                <ENTRY eventid="32" entrytime="00:01:04.19" heatid="32010" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2284" eventid="44" swimtime="00:00:29.38" lane="1" heatid="44014" points="323" />
                <RESULT resultid="2285" eventid="48" swimtime="00:01:09.00" lane="2" heatid="48003" points="343">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2286" eventid="52" status="DNS" swimtime="00:00:00.00" lane="3" heatid="52004" />
                <RESULT resultid="2287" eventid="32" swimtime="00:01:03.03" lane="2" heatid="32010" points="360">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2288" eventid="36" swimtime="00:02:29.65" lane="3" heatid="36002" points="351">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:54.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="496" birthdate="2010-01-01" gender="F" lastname="Frohlichová" firstname="Michaela" license="0" nation="GER">
              <ENTRIES>
                <ENTRY eventid="41" entrytime="00:00:32.29" heatid="41000" lane="0" />
                <ENTRY eventid="45" entrytime="00:01:28.68" heatid="45000" lane="0" />
                <ENTRY eventid="53" entrytime="00:02:41.70" heatid="53000" lane="0" />
                <ENTRY eventid="27" entrytime="00:00:41.17" heatid="27000" lane="0" />
                <ENTRY eventid="33" entrytime="00:01:16.24" heatid="33000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="2289" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="2290" eventid="33" status="WDR" swimtime="00:00:00.00" lane="0" heatid="33000" />
                <RESULT resultid="2291" eventid="41" status="WDR" swimtime="00:00:00.00" lane="0" heatid="41000" />
                <RESULT resultid="2292" eventid="45" status="WDR" swimtime="00:00:00.00" lane="0" heatid="45000" />
                <RESULT resultid="2293" eventid="53" status="WDR" swimtime="00:00:00.00" lane="0" heatid="53000" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:02:05.00" lane="1" heatid="11003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="849" eventid="11" swimtime="00:02:08.56" lane="1" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:04.25" />
                    <SPLIT distance="150" swimtime="00:01:38.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="245" number="1" />
                    <RELAYPOSITION athleteid="213" number="2" />
                    <RELAYPOSITION athleteid="253" number="3" />
                    <RELAYPOSITION athleteid="230" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="10" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:01:42.00" lane="1" heatid="40003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="850" eventid="40" status="DSQ" swimtime="00:01:38.75" lane="1" heatid="40003" comment="Die startenden Schwimmer, entsprechen nicht der im Meldeergebnis festgelegten Reihenfolge. Es nahmen nicht gemeldete Schwimmer teil.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.09" />
                    <SPLIT distance="100" swimtime="00:00:49.46" />
                    <SPLIT distance="150" swimtime="00:01:14.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="221" number="1" />
                    <RELAYPOSITION athleteid="220" number="2" />
                    <RELAYPOSITION athleteid="495" number="3" />
                    <RELAYPOSITION athleteid="258" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="11" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="71" entrytime="00:02:12.00" lane="1" heatid="71003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="851" eventid="71" swimtime="00:02:06.73" lane="1" heatid="71003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:39.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="254" number="1" />
                    <RELAYPOSITION athleteid="252" number="2" />
                    <RELAYPOSITION athleteid="259" number="3" />
                    <RELAYPOSITION athleteid="257" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="12" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="72" entrytime="00:01:51.10" lane="1" heatid="72003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="852" eventid="72" swimtime="00:01:48.02" lane="1" heatid="72003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.09" />
                    <SPLIT distance="100" swimtime="00:00:57.51" />
                    <SPLIT distance="150" swimtime="00:01:23.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="222" number="1" />
                    <RELAYPOSITION athleteid="256" number="2" />
                    <RELAYPOSITION athleteid="251" number="3" />
                    <RELAYPOSITION athleteid="260" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="13" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="72" entrytime="00:00:00.00" lane="1" heatid="72001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="853" eventid="72" swimtime="00:01:53.99" lane="1" heatid="72001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                    <SPLIT distance="100" swimtime="00:01:01.06" />
                    <SPLIT distance="150" swimtime="00:01:28.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="233" number="1" />
                    <RELAYPOSITION athleteid="221" number="2" />
                    <RELAYPOSITION athleteid="238" number="3" />
                    <RELAYPOSITION athleteid="255" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="14" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="72" entrytime="00:00:00.00" lane="4" heatid="72001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="854" eventid="72" swimtime="00:02:02.78" lane="4" heatid="72001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                    <SPLIT distance="150" swimtime="00:01:36.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="495" number="1" />
                    <RELAYPOSITION athleteid="220" number="2" />
                    <RELAYPOSITION athleteid="258" number="3" />
                    <RELAYPOSITION athleteid="226" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:00:00.00" lane="4" heatid="11001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="855" eventid="11" swimtime="00:02:35.48" lane="4" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                    <SPLIT distance="100" swimtime="00:01:14.58" />
                    <SPLIT distance="150" swimtime="00:01:55.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="250" number="1" />
                    <RELAYPOSITION athleteid="225" number="2" />
                    <RELAYPOSITION athleteid="231" number="3" />
                    <RELAYPOSITION athleteid="248" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:00:00.00" lane="1" heatid="11001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="856" eventid="11" swimtime="00:02:16.80" lane="1" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                    <SPLIT distance="150" swimtime="00:01:42.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="224" number="1" />
                    <RELAYPOSITION athleteid="237" number="2" />
                    <RELAYPOSITION athleteid="247" number="3" />
                    <RELAYPOSITION athleteid="261" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="23" entrytime="00:02:23.00" lane="4" heatid="23003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="857" eventid="23" status="DSQ" swimtime="00:02:28.76" lane="4" heatid="23003" comment="Beim Zielanschlag der Teilstrecke Brust hat der Sportler mit aufeinandergelegten Händen angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:01:57.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="213" number="1" />
                    <RELAYPOSITION athleteid="224" number="2" />
                    <RELAYPOSITION athleteid="253" number="3" />
                    <RELAYPOSITION athleteid="230" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="5" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="23" entrytime="00:00:00.00" lane="1" heatid="23001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="858" eventid="23" swimtime="00:02:34.56" lane="1" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="150" swimtime="00:01:59.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="219" number="1" />
                    <RELAYPOSITION athleteid="237" number="2" />
                    <RELAYPOSITION athleteid="245" number="3" />
                    <RELAYPOSITION athleteid="247" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="6" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="23" entrytime="00:00:00.00" lane="3" heatid="23001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="859" eventid="23" swimtime="00:02:47.45" lane="3" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:34.03" />
                    <SPLIT distance="150" swimtime="00:02:12.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="225" number="1" />
                    <RELAYPOSITION athleteid="242" number="2" />
                    <RELAYPOSITION athleteid="494" number="3" />
                    <RELAYPOSITION athleteid="261" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="7" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="39" entrytime="00:01:58.50" lane="1" heatid="39003" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="860" eventid="39" swimtime="00:01:53.87" lane="1" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:00:58.24" />
                    <SPLIT distance="150" swimtime="00:01:27.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="240" number="1" />
                    <RELAYPOSITION athleteid="254" number="2" />
                    <RELAYPOSITION athleteid="259" number="3" />
                    <RELAYPOSITION athleteid="257" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="8" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:00:00.00" lane="4" heatid="40001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="861" eventid="40" status="DSQ" swimtime="00:01:51.69" lane="4" heatid="40001" comment="Die startenden Schwimmer, entsprechen nicht der im Meldeergebnis festgelegten Reihenfolge. Es nahmen nicht gemeldete Schwimmer teil.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                    <SPLIT distance="100" swimtime="00:00:56.72" />
                    <SPLIT distance="150" swimtime="00:01:25.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="255" number="1" />
                    <RELAYPOSITION athleteid="251" number="2" />
                    <RELAYPOSITION athleteid="256" number="3" />
                    <RELAYPOSITION athleteid="260" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="9" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:00:00.00" lane="1" heatid="40001" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="862" eventid="40" swimtime="00:01:46.41" lane="1" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.68" />
                    <SPLIT distance="100" swimtime="00:00:52.82" />
                    <SPLIT distance="150" swimtime="00:01:19.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="222" number="1" />
                    <RELAYPOSITION athleteid="226" number="2" />
                    <RELAYPOSITION athleteid="233" number="3" />
                    <RELAYPOSITION athleteid="238" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSV Einheit Süd Chemnitz e.V." nation="GER" region="12" code="3403">
          <ATHLETES>
            <ATHLETE athleteid="347" birthdate="2015-01-01" gender="M" lastname="Barth" firstname="Romeo" license="484811" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:54.88" heatid="4003" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:44.36" heatid="8006" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:55.82" heatid="18004" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1556" eventid="4" swimtime="00:00:53.93" lane="4" heatid="4003" points="68" />
                <RESULT resultid="1557" eventid="8" swimtime="00:00:44.90" lane="4" heatid="8006" points="90" />
                <RESULT resultid="1558" eventid="18" status="DSQ" swimtime="00:00:55.77" lane="1" heatid="18004" comment="Beim Beinschlag wurden die Füße in der Rückwärtsbewegung nicht auswärts gedreht." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="348" birthdate="2011-01-01" gender="F" lastname="Friedrich" firstname="Laila" license="484803" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:35.03" heatid="43003" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:41.66" heatid="27007" lane="4" />
                <ENTRY eventid="33" entrytime="00:01:29.09" heatid="33003" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:41.23" heatid="41002" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:19.22" heatid="31003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1559" eventid="43" swimtime="00:00:34.92" lane="3" heatid="43003" points="283" />
                <RESULT resultid="1560" eventid="27" swimtime="00:00:41.85" lane="4" heatid="27007" points="311" />
                <RESULT resultid="1561" eventid="33" swimtime="00:01:29.75" lane="4" heatid="33003" points="249">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1562" eventid="41" swimtime="00:00:42.75" lane="1" heatid="41002" points="185" />
                <RESULT resultid="1563" eventid="31" swimtime="00:01:17.51" lane="4" heatid="31003" points="272">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="349" birthdate="2012-01-01" gender="M" lastname="Friedrich" firstname="Lenny" license="448794" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:41.82" heatid="4010" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:36.70" heatid="8013" lane="4" />
                <ENTRY eventid="18" entrytime="00:00:50.43" heatid="18006" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:24.67" heatid="20010" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1564" eventid="4" swimtime="00:00:42.43" lane="4" heatid="4010" points="141" />
                <RESULT resultid="1565" eventid="8" swimtime="00:00:38.58" lane="4" heatid="8013" points="142" />
                <RESULT resultid="1566" eventid="18" swimtime="00:00:55.87" lane="3" heatid="18006" points="89" />
                <RESULT resultid="1567" eventid="20" swimtime="00:01:27.15" lane="2" heatid="20010" points="136">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="350" birthdate="2013-01-01" gender="F" lastname="Graube" firstname="Freyja" license="484799" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:53.24" heatid="3007" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:40.73" heatid="7015" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:46.36" heatid="17014" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1568" eventid="3" swimtime="00:00:51.43" lane="2" heatid="3007" points="118" />
                <RESULT resultid="1569" eventid="7" swimtime="00:00:39.60" lane="3" heatid="7015" points="194" />
                <RESULT resultid="1570" eventid="17" swimtime="00:00:46.62" lane="3" heatid="17014" points="225" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="351" birthdate="2008-01-01" gender="F" lastname="Hänig" firstname="Lilly" license="428120">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:32.31" heatid="43005" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:40.48" heatid="27009" lane="1" />
                <ENTRY eventid="33" entrytime="00:01:26.43" heatid="33009" lane="4" />
                <ENTRY eventid="41" entrytime="00:00:39.04" heatid="41003" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:30.25" heatid="45007" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:17.42" heatid="31004" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1571" eventid="43" swimtime="00:00:33.02" lane="2" heatid="43005" points="334" />
                <RESULT resultid="1572" eventid="27" swimtime="00:00:41.91" lane="1" heatid="27009" points="310" />
                <RESULT resultid="1573" eventid="33" swimtime="00:01:28.25" lane="4" heatid="33009" points="262">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1574" eventid="41" swimtime="00:00:38.77" lane="2" heatid="41003" points="248" />
                <RESULT resultid="1575" eventid="45" swimtime="00:01:32.37" lane="4" heatid="45007" points="307">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1576" eventid="31" swimtime="00:01:17.00" lane="4" heatid="31004" points="277">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="352" birthdate="2015-01-01" gender="M" lastname="Karaus" firstname="Devin" license="484815" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:52.02" heatid="4003" lane="2" />
                <ENTRY eventid="6" entrytime="00:01:54.70" heatid="6003" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:39.74" heatid="8011" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1577" eventid="4" status="DNS" swimtime="00:00:00.00" lane="2" heatid="4003" />
                <RESULT resultid="1578" eventid="6" status="DNS" swimtime="00:00:00.00" lane="1" heatid="6003" />
                <RESULT resultid="1579" eventid="8" status="DNS" swimtime="00:00:00.00" lane="4" heatid="8011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="353" birthdate="2012-01-01" gender="M" lastname="Karaus" firstname="Lenjo" license="448793" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:43.77" heatid="4009" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:35.21" heatid="8014" lane="2" />
                <ENTRY eventid="10" entrytime="00:01:31.78" heatid="10005" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1580" eventid="4" status="DNS" swimtime="00:00:00.00" lane="4" heatid="4009" />
                <RESULT resultid="1581" eventid="8" status="DNS" swimtime="00:00:00.00" lane="2" heatid="8014" />
                <RESULT resultid="1582" eventid="10" status="DNS" swimtime="00:00:00.00" lane="3" heatid="10005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="354" birthdate="2013-01-01" gender="M" lastname="Klötzner" firstname="Jaden Pascal" license="471866" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:49.77" heatid="4005" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:38.83" heatid="8011" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:51.67" heatid="18006" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:32.08" heatid="20008" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1583" eventid="4" swimtime="00:00:51.84" lane="2" heatid="4005" points="77" />
                <RESULT resultid="1584" eventid="8" swimtime="00:00:40.81" lane="2" heatid="8011" points="120" />
                <RESULT resultid="1585" eventid="18" swimtime="00:00:55.37" lane="1" heatid="18006" points="91" />
                <RESULT resultid="1586" eventid="20" swimtime="00:01:33.40" lane="4" heatid="20008" points="110">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="355" birthdate="2006-01-01" gender="F" lastname="Köhler" firstname="Lea Sophie" license="387692">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:30.11" heatid="43014" lane="1" />
                <ENTRY eventid="33" entrytime="00:01:16.48" heatid="33010" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:32.08" heatid="41012" lane="1" />
                <ENTRY eventid="45" entrytime="00:01:26.14" heatid="45008" lane="3" />
                <ENTRY eventid="53" entrytime="00:02:54.79" heatid="53001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1587" eventid="43" swimtime="00:00:30.97" lane="1" heatid="43014" points="405" />
                <RESULT resultid="1588" eventid="33" swimtime="00:01:19.09" lane="1" heatid="33010" points="364">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1589" eventid="41" swimtime="00:00:32.91" lane="1" heatid="41012" points="406" />
                <RESULT resultid="1590" eventid="45" swimtime="00:01:26.38" lane="3" heatid="45008" points="376">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1591" eventid="53" swimtime="00:03:05.97" lane="2" heatid="53001" points="281">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.60" />
                    <SPLIT distance="100" swimtime="00:01:27.61" />
                    <SPLIT distance="150" swimtime="00:02:19.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="356" birthdate="1992-01-01" gender="M" lastname="Metzner" firstname="Joshua" license="149240">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:25.13" heatid="44013" lane="4" />
                <ENTRY eventid="48" entrytime="00:01:03.25" heatid="48006" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:27.36" heatid="42008" lane="1" />
                <ENTRY eventid="26" entrytime="00:00:29.67" heatid="26005" lane="3" />
                <ENTRY eventid="36" entrytime="00:02:21.12" heatid="36003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1592" eventid="44" swimtime="00:00:26.09" lane="4" heatid="44013" points="461" />
                <RESULT resultid="1593" eventid="48" swimtime="00:01:03.86" lane="2" heatid="48006" points="433">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1594" eventid="42" swimtime="00:00:27.30" lane="1" heatid="42008" points="505" />
                <RESULT resultid="1595" eventid="26" swimtime="00:00:29.75" lane="3" heatid="26005" points="410" />
                <RESULT resultid="1596" eventid="36" swimtime="00:02:24.38" lane="4" heatid="36003" points="391">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:09.15" />
                    <SPLIT distance="150" swimtime="00:01:46.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="357" birthdate="2009-01-01" gender="F" lastname="Rudolph" firstname="Anna" license="386529">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:34.23" heatid="43004" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:43.04" heatid="27004" lane="1" />
                <ENTRY eventid="33" entrytime="00:01:29.33" heatid="33002" lane="2" />
                <ENTRY eventid="45" entrytime="00:01:33.84" heatid="45003" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:17.28" heatid="31004" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1597" eventid="43" swimtime="00:00:35.15" lane="3" heatid="43004" points="277" />
                <RESULT resultid="1598" eventid="27" swimtime="00:00:43.74" lane="1" heatid="27004" points="272" />
                <RESULT resultid="1599" eventid="33" swimtime="00:01:31.57" lane="2" heatid="33002" points="235">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1600" eventid="45" swimtime="00:01:36.02" lane="3" heatid="45003" points="273">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1601" eventid="31" swimtime="00:01:19.02" lane="1" heatid="31004" points="257">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="358" birthdate="2013-01-01" gender="M" lastname="Schönberg" firstname="Noah" license="453239" nation="GER" easy.nation2="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:43.75" heatid="4009" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:36.87" heatid="8012" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:46.99" heatid="18007" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:25.96" heatid="20010" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1602" eventid="4" swimtime="00:00:43.69" lane="1" heatid="4009" points="129" />
                <RESULT resultid="1603" eventid="8" swimtime="00:00:36.69" lane="2" heatid="8012" points="165" />
                <RESULT resultid="1604" eventid="18" swimtime="00:00:48.46" lane="1" heatid="18007" points="136" />
                <RESULT resultid="1605" eventid="20" swimtime="00:01:24.69" lane="4" heatid="20010" points="148">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="359" birthdate="2010-01-01" gender="M" lastname="Schulz" firstname="John" license="448791" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:33.15" heatid="44003" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:47.01" heatid="28001" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:39.78" heatid="42001" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:41.65" heatid="26001" lane="2" />
                <ENTRY eventid="32" entrytime="00:01:14.77" heatid="32002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1606" eventid="44" swimtime="00:00:32.67" lane="4" heatid="44003" points="234" />
                <RESULT resultid="1607" eventid="28" swimtime="00:00:44.62" lane="1" heatid="28001" points="174" />
                <RESULT resultid="1608" eventid="42" swimtime="00:00:39.85" lane="2" heatid="42001" points="162" />
                <RESULT resultid="1609" eventid="26" swimtime="00:00:40.64" lane="2" heatid="26001" points="161" />
                <RESULT resultid="1610" eventid="32" swimtime="00:01:14.96" lane="3" heatid="32002" points="214">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="360" birthdate="2011-01-01" gender="M" lastname="Spielvogel" firstname="Oskar" license="449485" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:36.82" heatid="44001" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:49.17" heatid="28001" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:41.68" heatid="42001" lane="3" />
                <ENTRY eventid="26" entrytime="00:00:52.11" heatid="26001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1611" eventid="44" swimtime="00:00:36.09" lane="3" heatid="44001" points="174" />
                <RESULT resultid="1612" eventid="28" swimtime="00:00:49.66" lane="4" heatid="28001" points="126" />
                <RESULT resultid="1613" eventid="42" swimtime="00:00:43.57" lane="3" heatid="42001" points="124" />
                <RESULT resultid="1614" eventid="26" swimtime="00:00:45.86" lane="1" heatid="26001" points="112" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Ústecká akademie plaveckých sportu z.s." nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="185" birthdate="2007-01-01" gender="M" lastname="Adamec" firstname="Petr" license="38760000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.26" heatid="44000" lane="0" />
                <ENTRY eventid="52" entrytime="00:01:55.21" heatid="52000" lane="0" />
                <ENTRY eventid="32" entrytime="00:00:52.43" heatid="32000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="834" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="835" eventid="52" status="WDR" swimtime="00:00:00.00" lane="0" heatid="52000" />
                <RESULT resultid="836" eventid="32" status="WDR" swimtime="00:00:00.00" lane="0" heatid="32000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="186" birthdate="2008-01-01" gender="M" lastname="Bartuska" firstname="Daniel" license="42309000">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:32.91" heatid="28010" lane="1" />
                <ENTRY eventid="30" entrytime="00:01:09.04" heatid="30005" lane="4" />
                <ENTRY eventid="38" entrytime="00:02:37.16" heatid="38005" lane="3" />
                <ENTRY eventid="42" entrytime="00:00:29.02" heatid="42006" lane="1" />
                <ENTRY eventid="46" entrytime="00:01:11.21" heatid="46006" lane="1" />
                <ENTRY eventid="54" entrytime="00:02:21.86" heatid="54004" lane="3" />
                <ENTRY eventid="61" entrytime="00:00:32.46" heatid="61001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="837" eventid="28" swimtime="00:00:32.46" lane="1" heatid="28010" points="454" />
                <RESULT resultid="838" eventid="30" swimtime="00:01:05.93" lane="4" heatid="30005" points="380">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="839" eventid="38" swimtime="00:02:36.73" lane="3" heatid="38005" points="450">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="150" swimtime="00:01:56.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="840" eventid="42" swimtime="00:00:28.03" lane="1" heatid="42006" points="467" />
                <RESULT resultid="841" eventid="46" swimtime="00:01:11.42" lane="1" heatid="46006" points="463">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="842" eventid="54" swimtime="00:02:24.38" lane="3" heatid="54004" points="437">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:10.19" />
                    <SPLIT distance="150" swimtime="00:01:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2326" eventid="61" swimtime="00:00:32.61" lane="4" heatid="61001" points="447" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="187" birthdate="2004-01-01" gender="M" lastname="Beca" firstname="Jakub" license="35985000">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:24.17" heatid="44017" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:31.57" heatid="28007" lane="2" />
                <ENTRY eventid="42" entrytime="00:00:25.89" heatid="42009" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:26.35" heatid="26010" lane="3" />
                <ENTRY eventid="58" entrytime="00:00:26.60" heatid="58001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="843" eventid="44" swimtime="00:00:24.22" lane="4" heatid="44017" points="576" />
                <RESULT resultid="844" eventid="28" swimtime="00:00:31.50" lane="2" heatid="28007" points="496" />
                <RESULT resultid="845" eventid="42" swimtime="00:00:25.79" lane="2" heatid="42009" points="599" />
                <RESULT resultid="846" eventid="26" swimtime="00:00:26.60" lane="3" heatid="26010" points="574" />
                <RESULT resultid="2360" eventid="58" swimtime="00:00:26.35" lane="3" heatid="58001" points="590" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="188" birthdate="1999-01-01" gender="F" lastname="Plihalova" firstname="Anna" license="25260000">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:31.75" heatid="27009" lane="4" />
                <ENTRY eventid="45" entrytime="00:01:09.64" heatid="45008" lane="2" />
                <ENTRY eventid="60" entrytime="00:00:32.06" heatid="60001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="847" eventid="27" swimtime="00:00:32.06" lane="4" heatid="27009" points="692" />
                <RESULT resultid="848" eventid="45" swimtime="00:01:09.21" lane="2" heatid="45008" points="731">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2319" eventid="60" swimtime="00:00:31.51" lane="2" heatid="60001" points="729" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="WSG Jena-Lobeda e.V." nation="GER" region="16" code="3278">
          <ATHLETES>
            <ATHLETE athleteid="14" birthdate="2012-01-01" gender="F" lastname="Brose" firstname="Frieda Barbara" license="505004" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:37.46" heatid="43002" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:39.35" heatid="27006" lane="2" />
                <ENTRY eventid="37" entrytime="00:03:15.72" heatid="37001" lane="3" />
                <ENTRY eventid="45" entrytime="00:01:29.06" heatid="45004" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="57" eventid="43" swimtime="00:00:36.19" lane="1" heatid="43002" points="254" />
                <RESULT resultid="58" eventid="27" swimtime="00:00:39.73" lane="2" heatid="27006" points="364" />
                <RESULT resultid="59" eventid="37" swimtime="00:03:10.14" lane="3" heatid="37001" points="354">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                    <SPLIT distance="100" swimtime="00:01:33.45" />
                    <SPLIT distance="150" swimtime="00:02:23.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="60" eventid="45" swimtime="00:01:29.80" lane="3" heatid="45004" points="334">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="15" birthdate="2010-01-01" gender="M" lastname="Chegrakhcy" firstname="Serhii" license="491079" nation="UKR">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:27.44" heatid="44009" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:30.08" heatid="42005" lane="1" />
                <ENTRY eventid="32" entrytime="00:01:00.39" heatid="32007" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="61" eventid="44" swimtime="00:00:27.36" lane="1" heatid="44009" points="400" />
                <RESULT resultid="62" eventid="42" swimtime="00:00:30.14" lane="1" heatid="42005" points="375" />
                <RESULT resultid="63" eventid="32" swimtime="00:01:01.41" lane="3" heatid="32007" points="389">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="16" birthdate="2012-01-01" gender="F" lastname="Greinke" firstname="Magdalena Ruth" license="458790" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:37.90" heatid="43001" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:49.24" heatid="27001" lane="4" />
                <ENTRY eventid="25" entrytime="00:00:45.62" heatid="25001" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:27.53" heatid="31001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="64" eventid="43" swimtime="00:00:36.56" lane="1" heatid="43001" points="246" />
                <RESULT resultid="65" eventid="27" swimtime="00:00:47.83" lane="4" heatid="27001" points="208" />
                <RESULT resultid="66" eventid="25" swimtime="00:00:43.67" lane="1" heatid="25001" points="193" />
                <RESULT resultid="67" eventid="31" swimtime="00:01:27.16" lane="3" heatid="31001" points="191">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="17" birthdate="2010-01-01" gender="F" lastname="Grimmer" firstname="Rita" license="446916" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:32.74" heatid="43000" lane="0" />
                <ENTRY eventid="33" entrytime="00:01:30.62" heatid="33000" lane="0" />
                <ENTRY eventid="31" entrytime="00:01:17.33" heatid="31000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="68" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
                <RESULT resultid="69" eventid="33" status="WDR" swimtime="00:00:00.00" lane="0" heatid="33000" />
                <RESULT resultid="70" eventid="31" status="WDR" swimtime="00:00:00.00" lane="0" heatid="31000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="18" birthdate="1995-01-01" gender="F" lastname="Kammel" firstname="Sarah" license="169382" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:32.16" heatid="43014" lane="4" />
                <ENTRY eventid="25" entrytime="00:00:38.18" heatid="25009" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:13.31" heatid="31013" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="71" eventid="43" status="WDR" swimtime="00:00:00.00" lane="4" heatid="43014" />
                <RESULT resultid="72" eventid="25" status="WDR" swimtime="00:00:00.00" lane="1" heatid="25009" />
                <RESULT resultid="73" eventid="31" status="WDR" swimtime="00:00:00.00" lane="4" heatid="31013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="19" birthdate="2013-01-01" gender="M" lastname="Kochzius" firstname="Albert" license="458791" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:41.44" heatid="6011" lane="4" />
                <ENTRY eventid="16" entrytime="00:01:30.96" heatid="16010" lane="1" />
                <ENTRY eventid="18" entrytime="00:00:44.06" heatid="18014" lane="4" />
                <ENTRY eventid="38" entrytime="00:03:35.14" heatid="38002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="74" eventid="6" swimtime="00:01:41.53" lane="4" heatid="6011" points="161">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="75" eventid="16" swimtime="00:01:30.57" lane="1" heatid="16010" points="151">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="76" eventid="18" swimtime="00:00:46.74" lane="4" heatid="18014" points="152" />
                <RESULT resultid="77" eventid="38" swimtime="00:03:29.65" lane="2" heatid="38002" points="188">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.15" />
                    <SPLIT distance="100" swimtime="00:01:40.49" />
                    <SPLIT distance="150" swimtime="00:02:34.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="20" birthdate="2014-01-01" gender="F" lastname="Kölling" firstname="Lisa" license="464910" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:39.84" heatid="5010" lane="4" />
                <ENTRY eventid="9" entrytime="00:01:34.44" heatid="9010" lane="3" />
                <ENTRY eventid="17" entrytime="00:00:45.43" heatid="17015" lane="4" />
                <ENTRY eventid="37" entrytime="00:03:39.07" heatid="37001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="78" eventid="5" swimtime="00:01:38.95" lane="4" heatid="5010" points="250">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="79" eventid="9" swimtime="00:01:35.31" lane="3" heatid="9010" points="208">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="80" eventid="17" swimtime="00:00:45.49" lane="4" heatid="17015" points="242" />
                <RESULT resultid="81" eventid="37" swimtime="00:03:30.20" lane="4" heatid="37001" points="262">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                    <SPLIT distance="100" swimtime="00:01:42.79" />
                    <SPLIT distance="150" swimtime="00:02:37.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="21" birthdate="2010-01-01" gender="M" lastname="Kovezin" firstname="Vladimir" license="423550" nation="GER">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:39.65" heatid="28004" lane="4" />
                <ENTRY eventid="34" entrytime="00:01:19.94" heatid="34003" lane="3" />
                <ENTRY eventid="46" entrytime="00:01:25.83" heatid="46002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="82" eventid="28" swimtime="00:00:38.42" lane="4" heatid="28004" points="273" />
                <RESULT resultid="83" eventid="34" swimtime="00:01:19.12" lane="3" heatid="34003" points="241">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="84" eventid="46" swimtime="00:01:27.65" lane="4" heatid="46002" points="250">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="22" birthdate="2008-01-01" gender="M" lastname="Lindemann" firstname="Aron" license="393036" nation="GER">
              <ENTRIES>
                <ENTRY eventid="28" entrytime="00:00:34.65" heatid="28005" lane="3" />
                <ENTRY eventid="34" entrytime="00:01:10.28" heatid="34008" lane="4" />
                <ENTRY eventid="46" entrytime="00:01:17.70" heatid="46002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="85" eventid="28" swimtime="00:00:33.83" lane="3" heatid="28005" points="401" />
                <RESULT resultid="86" eventid="34" swimtime="00:01:11.26" lane="4" heatid="34008" points="330">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="87" eventid="46" swimtime="00:01:15.66" lane="2" heatid="46002" points="390">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="23" birthdate="2007-01-01" gender="F" lastname="Lippert" firstname="Josephine" license="383842" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:33.74" heatid="43004" lane="2" />
                <ENTRY eventid="47" entrytime="00:01:26.82" heatid="47007" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:17.48" heatid="31003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="88" eventid="43" status="WDR" swimtime="00:00:00.00" lane="2" heatid="43004" />
                <RESULT resultid="89" eventid="47" status="WDR" swimtime="00:00:00.00" lane="4" heatid="47007" />
                <RESULT resultid="90" eventid="31" status="WDR" swimtime="00:00:00.00" lane="2" heatid="31003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="24" birthdate="2012-01-01" gender="M" lastname="Lorenz" firstname="Theo" license="458792" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:39.09" heatid="4016" lane="2" />
                <ENTRY eventid="8" entrytime="00:00:36.33" heatid="8013" lane="3" />
                <ENTRY eventid="16" entrytime="00:01:27.27" heatid="16011" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:24.42" heatid="20011" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="91" eventid="4" swimtime="00:00:36.28" lane="2" heatid="4016" points="226" />
                <RESULT resultid="92" eventid="8" swimtime="00:00:34.79" lane="3" heatid="8013" points="194" />
                <RESULT resultid="93" eventid="16" swimtime="00:01:23.95" lane="3" heatid="16011" points="190">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="94" eventid="20" swimtime="00:01:18.98" lane="4" heatid="20011" points="182">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="25" birthdate="2014-01-01" gender="F" lastname="Meierkord" firstname="Rachel" license="468845" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:37.63" heatid="5010" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:34.51" heatid="9010" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:44.36" heatid="17015" lane="2" />
                <ENTRY eventid="37" entrytime="00:03:30.76" heatid="37001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="95" eventid="5" swimtime="00:01:36.63" lane="1" heatid="5010" points="268">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="96" eventid="9" swimtime="00:01:31.34" lane="1" heatid="9010" points="236">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="97" eventid="17" swimtime="00:00:44.40" lane="2" heatid="17015" points="260" />
                <RESULT resultid="98" eventid="37" swimtime="00:03:28.47" lane="1" heatid="37001" points="268">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:42.44" />
                    <SPLIT distance="150" swimtime="00:02:36.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="26" birthdate="2011-01-01" gender="F" lastname="Mutschke" firstname="Luisa" license="442362" nation="GER">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:46.81" heatid="27001" lane="2" />
                <ENTRY eventid="33" entrytime="00:01:29.03" heatid="33003" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:18.30" heatid="31003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="99" eventid="27" swimtime="00:00:47.24" lane="2" heatid="27001" points="216" />
                <RESULT resultid="100" eventid="33" status="DSQ" swimtime="00:01:30.73" lane="1" heatid="33003" comment="Die Teilstrecke Rücken wurde nicht in Rückenlage beendet.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="101" eventid="31" swimtime="00:01:18.98" lane="3" heatid="31003" points="257">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="27" birthdate="2013-01-01" gender="F" lastname="Mutschke" firstname="Sarah" license="464904" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:45.26" heatid="5008" lane="4" />
                <ENTRY eventid="7" entrytime="00:00:38.16" heatid="7018" lane="1" />
                <ENTRY eventid="17" entrytime="00:00:47.43" heatid="17013" lane="3" />
                <ENTRY eventid="19" entrytime="00:01:34.26" heatid="19011" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="102" eventid="5" swimtime="00:01:42.88" lane="4" heatid="5008" points="222">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="103" eventid="7" swimtime="00:00:36.39" lane="1" heatid="7018" points="250" />
                <RESULT resultid="104" eventid="17" swimtime="00:00:45.27" lane="3" heatid="17013" points="246" />
                <RESULT resultid="105" eventid="19" swimtime="00:01:28.71" lane="2" heatid="19011" points="181">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="28" birthdate="2009-01-01" gender="M" lastname="Neuhaus" firstname="Jakob Friedrich" license="437045" nation="GER">
              <ENTRIES>
                <ENTRY eventid="30" entrytime="00:01:15.19" heatid="30001" lane="3" />
                <ENTRY eventid="34" entrytime="00:01:16.92" heatid="34004" lane="1" />
                <ENTRY eventid="26" entrytime="00:00:38.52" heatid="26002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="106" eventid="30" swimtime="00:01:15.12" lane="3" heatid="30001" points="257">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="107" eventid="34" swimtime="00:01:17.54" lane="1" heatid="34004" points="256">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="108" eventid="26" swimtime="00:00:34.90" lane="1" heatid="26002" points="254" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="29" birthdate="2014-01-01" gender="F" lastname="Raymundo" firstname="Emilia Katerina" license="458887" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:33.91" heatid="5014" lane="1" />
                <ENTRY eventid="9" entrytime="00:01:22.90" heatid="9017" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:14.82" heatid="19020" lane="2" />
                <ENTRY eventid="21" entrytime="00:03:04.16" heatid="21004" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="109" eventid="5" swimtime="00:01:31.34" lane="1" heatid="5014" points="318">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="110" eventid="9" swimtime="00:01:20.04" lane="2" heatid="9017" points="351">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="111" eventid="19" swimtime="00:01:13.58" lane="2" heatid="19020" points="318">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="112" eventid="21" swimtime="00:02:58.59" lane="1" heatid="21004" points="317">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:22.73" />
                    <SPLIT distance="150" swimtime="00:02:15.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="30" birthdate="2013-01-01" gender="M" lastname="Schmidt" firstname="Robert" license="458795" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:23.24" heatid="2005" lane="1" />
                <ENTRY eventid="8" entrytime="00:00:30.11" heatid="8024" lane="1" />
                <ENTRY eventid="20" entrytime="00:01:10.34" heatid="20021" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="113" eventid="2" swimtime="00:01:21.26" lane="1" heatid="2005" points="203">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="114" eventid="8" swimtime="00:00:29.64" lane="1" heatid="8024" points="314" />
                <RESULT resultid="115" eventid="20" swimtime="00:01:09.53" lane="1" heatid="20021" points="268">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="31" birthdate="2014-01-01" gender="F" lastname="Schönfeld" firstname="Viola" license="464905" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:52.92" heatid="5005" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:35.83" heatid="7023" lane="4" />
                <ENTRY eventid="17" entrytime="00:00:45.43" heatid="17015" lane="1" />
                <ENTRY eventid="19" entrytime="00:01:23.79" heatid="19016" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="116" eventid="5" swimtime="00:01:36.56" lane="2" heatid="5005" points="269">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="117" eventid="7" swimtime="00:00:34.42" lane="4" heatid="7023" points="295" />
                <RESULT resultid="118" eventid="17" swimtime="00:00:44.62" lane="1" heatid="17015" points="257" />
                <RESULT resultid="119" eventid="19" swimtime="00:01:19.78" lane="2" heatid="19016" points="249">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="32" birthdate="2011-01-01" gender="M" lastname="Simon" firstname="Bruno" license="442369" nation="GER">
              <ENTRIES>
                <ENTRY eventid="44" entrytime="00:00:39.20" heatid="44001" lane="1" />
                <ENTRY eventid="34" entrytime="00:01:25.26" heatid="34001" lane="2" />
                <ENTRY eventid="32" entrytime="00:01:17.27" heatid="32001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="120" eventid="44" swimtime="00:00:31.86" lane="1" heatid="44001" points="253" />
                <RESULT resultid="121" eventid="34" swimtime="00:01:23.21" lane="2" heatid="34001" points="207">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="122" eventid="32" swimtime="00:01:14.41" lane="2" heatid="32001" points="218">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="33" birthdate="2011-01-01" gender="F" lastname="Steiniger" firstname="Enne Therese" license="442367" nation="GER">
              <ENTRIES>
                <ENTRY eventid="43" entrytime="00:00:31.70" heatid="43006" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:25.08" heatid="47005" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:13.14" heatid="31010" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="123" eventid="43" swimtime="00:00:31.94" lane="3" heatid="43006" points="370" />
                <RESULT resultid="124" eventid="47" swimtime="00:01:24.29" lane="1" heatid="47005" points="276">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="125" eventid="31" swimtime="00:01:12.98" lane="4" heatid="31010" points="326">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="34" birthdate="2002-01-01" gender="F" lastname="Vorberger" firstname="Aina" license="290604" nation="GER">
              <ENTRIES>
                <ENTRY eventid="33" entrytime="00:01:13.57" heatid="33010" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:31.21" heatid="41012" lane="3" />
                <ENTRY eventid="49" entrytime="00:02:39.76" heatid="49001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="126" eventid="33" swimtime="00:01:15.25" lane="2" heatid="33010" points="423">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="127" eventid="41" swimtime="00:00:31.98" lane="3" heatid="41012" points="443" />
                <RESULT resultid="128" eventid="49" swimtime="00:02:50.70" lane="3" heatid="49001" points="344">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="150" swimtime="00:02:04.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="35" birthdate="2011-01-01" gender="F" lastname="Weber" firstname="Stella" license="462719" nation="GER">
              <ENTRIES>
                <ENTRY eventid="27" entrytime="00:00:44.13" heatid="27003" lane="1" />
                <ENTRY eventid="41" entrytime="00:00:38.52" heatid="41004" lane="1" />
                <ENTRY eventid="45" entrytime="00:01:35.01" heatid="45003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="129" eventid="27" status="WDR" swimtime="00:00:00.00" lane="1" heatid="27003" />
                <RESULT resultid="130" eventid="41" status="WDR" swimtime="00:00:00.00" lane="1" heatid="41004" />
                <RESULT resultid="131" eventid="45" status="WDR" swimtime="00:00:00.00" lane="1" heatid="45003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="ZKP Frankenstein Zabkowice Slaskie" nation="POL" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="361" birthdate="2012-01-01" gender="M" lastname="Antonyshyn" firstname="Maksym" license="0">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:00:46.90" heatid="8004" lane="2" />
                <ENTRY eventid="18" entrytime="00:00:52.30" heatid="18006" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1615" eventid="8" swimtime="00:00:40.25" lane="2" heatid="8004" points="125" />
                <RESULT resultid="1616" eventid="18" status="DNS" swimtime="00:00:00.00" lane="4" heatid="18006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="362" birthdate="2014-01-01" gender="M" lastname="Cyganek" firstname="Hubert" license="0">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:50.00" heatid="4005" lane="3" />
                <ENTRY eventid="8" entrytime="00:00:46.70" heatid="8005" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1617" eventid="4" status="DSQ" swimtime="00:00:54.84" lane="3" heatid="4005" comment="Der Sportler hat bei der Rückenstarthilfe nicht mit mind. einer Zehe jeden Fußes die Wand berührt." />
                <RESULT resultid="1618" eventid="8" swimtime="00:00:49.61" lane="1" heatid="8005" points="67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="363" birthdate="2012-01-01" gender="M" lastname="Cyganek" firstname="Julian" license="0">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:47.90" heatid="6004" lane="3" />
                <ENTRY eventid="18" entrytime="00:00:54.00" heatid="18005" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1619" eventid="6" swimtime="00:02:12.53" lane="3" heatid="6004" points="72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1620" eventid="18" status="DSQ" swimtime="00:00:57.60" lane="4" heatid="18005" comment="Beim Zielanschlag hat der Sportler nicht mit beiden Händen gleichzeitig angeschlagen." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="364" birthdate="2015-01-01" gender="F" lastname="Garbowska" firstname="Julia" license="0">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:00:54.00" heatid="3006" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:50.00" heatid="7007" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1621" eventid="3" status="DSQ" swimtime="00:01:05.29" lane="3" heatid="3006" comment="Die Sportlerin hat bei der  Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt." />
                <RESULT resultid="1622" eventid="7" status="DSQ" swimtime="00:01:03.33" lane="3" heatid="7007" comment="Die Sportlerin startete vor dem Startsignal" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="365" birthdate="2014-01-01" gender="M" lastname="Goryl" firstname="Aleksander" license="0">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:00:42.80" heatid="8007" lane="2" />
                <ENTRY eventid="14" entrytime="00:00:49.00" heatid="14003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1623" eventid="8" swimtime="00:00:42.99" lane="2" heatid="8007" points="103" />
                <RESULT resultid="1624" eventid="14" status="DSQ" swimtime="00:00:58.83" lane="1" heatid="14003" comment="Beim Anschlag an der Wende hat der Sportler nicht mit beiden Händen gleichzeitig angeschlagen." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="366" birthdate="2016-01-01" gender="F" lastname="Mackiewicz" firstname="Pola" license="0">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:00:47.20" heatid="7009" lane="2" />
                <ENTRY eventid="17" entrytime="00:00:51.20" heatid="17017" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1625" eventid="7" status="DNS" swimtime="00:00:00.00" lane="2" heatid="7009" />
                <RESULT resultid="1626" eventid="17" status="DNS" swimtime="00:00:00.00" lane="4" heatid="17017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="367" birthdate="2014-01-01" gender="M" lastname="Maj" firstname="Piotr" license="0">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:00:44.10" heatid="8006" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:34.50" heatid="20007" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1627" eventid="8" swimtime="00:00:37.31" lane="3" heatid="8006" points="157" />
                <RESULT resultid="1628" eventid="20" status="DSQ" swimtime="00:01:41.09" lane="3" heatid="20007" comment="Der Sportler startete vor dem Startsignal">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="368" birthdate="2017-01-01" gender="M" lastname="Malecki" firstname="Oskar" license="0">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:00:41.00" heatid="8020" lane="2" />
                <ENTRY eventid="20" entrytime="00:01:33.00" heatid="20017" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1629" eventid="8" status="DSQ" swimtime="00:00:40.91" lane="2" heatid="8020" comment="Der Sportler startete vor dem Startsignal" />
                <RESULT resultid="1630" eventid="20" swimtime="00:01:34.83" lane="2" heatid="20017" points="105">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="369" birthdate="2014-01-01" gender="M" lastname="Szczepaniak" firstname="Marcin" license="0">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:00:43.10" heatid="8007" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:34.70" heatid="20007" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1631" eventid="8" swimtime="00:00:42.34" lane="3" heatid="8007" points="107" />
                <RESULT resultid="1632" eventid="20" swimtime="00:01:40.54" lane="1" heatid="20007" points="88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST name="Pflichtzeiten 2015 weiblich" course="SCM" gender="F" timestandardlistid="1">
      <AGEGROUP agemax="10" agemin="10" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2014 weiblich" course="SCM" gender="F" timestandardlistid="2">
      <AGEGROUP agemax="11" agemin="11" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2013 weiblich" course="SCM" gender="F" timestandardlistid="3">
      <AGEGROUP agemax="12" agemin="12" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:34.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2015 männlich" course="SCM" gender="M" timestandardlistid="4">
      <AGEGROUP agemax="10" agemin="10" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2014 männlich" course="SCM" gender="M" timestandardlistid="5">
      <AGEGROUP agemax="11" agemin="11" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2013 männlich" course="SCM" gender="M" timestandardlistid="6">
      <AGEGROUP agemax="12" agemin="12" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:34.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2012 männlich" course="SCM" gender="M" timestandardlistid="7">
      <AGEGROUP agemax="13" agemin="13" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2017 weiblich" course="SCM" gender="F" timestandardlistid="8">
      <AGEGROUP agemax="8" agemin="8" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2016 weiblich" course="SCM" gender="F" timestandardlistid="9">
      <AGEGROUP agemax="9" agemin="9" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2017 männlich" course="SCM" gender="M" timestandardlistid="10">
      <AGEGROUP agemax="8" agemin="8" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2016 männlich" course="SCM" gender="M" timestandardlistid="11">
      <AGEGROUP agemax="9" agemin="9" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2006 und jünger männlich" course="SCM" gender="M" timestandardlistid="12">
      <AGEGROUP agemax="-1" agemin="19" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:18.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:18.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:16.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2011 männlich" course="SCM" gender="M" timestandardlistid="13">
      <AGEGROUP agemax="14" agemin="14" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:33.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:28.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2009 bis 2010 männlich" course="SCM" gender="M" timestandardlistid="14">
      <AGEGROUP agemax="16" agemin="15" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:26.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:24.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2007 bis 2008 männlich" course="SCM" gender="M" timestandardlistid="15">
      <AGEGROUP agemax="18" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:24.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2012 weiblich" course="SCM" gender="F" timestandardlistid="16">
      <AGEGROUP agemax="13" agemin="13" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2011 weiblich" course="SCM" gender="F" timestandardlistid="17">
      <AGEGROUP agemax="14" agemin="14" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:33.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:28.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:33.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:33.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:38.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2009 bis 2010 weiblich" course="SCM" gender="F" timestandardlistid="18">
      <AGEGROUP agemax="16" agemin="15" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:31.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:26.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:31.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:31.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:36.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2007 bis 2008 weiblich" course="SCM" gender="F" timestandardlistid="19">
      <AGEGROUP agemax="18" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:24.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2006 und jünger weiblich" course="SCM" gender="F" timestandardlistid="20">
      <AGEGROUP agemax="-1" agemin="19" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
