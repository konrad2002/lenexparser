<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.30" registration="Oliver Busch">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Halle (Saale)" course="LCM" name="Mitteldeutsche Meisterschaften" nation="GER" organizer="SV Halle e. V. Abteilung Schwimmen" hostclub="Landesschwimmverband Sachsen-Anhalt e. V." deadline="2025-06-23" timing="AUTOMATIC">
      <CONTACT email="ollibusch@freenet.de" name="Busch, Oliver" phone="0176 24840175" />
      <AGEDATE type="YEAR" value="2025-01-01" />
      <BANK name="Volksbank Halle/S. e. G." iban="DE37 8009 3784 0002 1234 52" bic="" accountholder="Landesschwimmverband Sachsen-Anhalt e. V." note="Mdt. Meisterschaften 2025 + Vereinsname" />
      <SESSIONS>
        <SESSION number="1" date="2025-07-05" daytime="10:00" officialmeeting="09:30" warmupfrom="08:30">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="F" round="PRE" order="1">
              <SWIMSTYLE name="100m Schmetterling weiblich (Vorlauf)" stroke="FLY" relaycount="1" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="1001" number="1" daytime="10:00" />
                <HEAT heatid="1002" number="2" daytime="10:02" />
                <HEAT heatid="1003" number="3" daytime="10:04" />
                <HEAT heatid="1004" number="4" daytime="10:06" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="688" />
                    <RANKING place="2" resultid="704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="196" />
                    <RANKING place="5" resultid="507" />
                    <RANKING place="4" resultid="612" />
                    <RANKING place="3" resultid="653" />
                    <RANKING place="2" resultid="773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="6" resultid="49" />
                    <RANKING place="5" resultid="153" />
                    <RANKING place="2" resultid="334" />
                    <RANKING place="3" resultid="396" />
                    <RANKING place="4" resultid="476" />
                    <RANKING place="7" resultid="584" />
                    <RANKING place="8" resultid="607" />
                    <RANKING place="1" resultid="618" />
                    <RANKING place="9" resultid="625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="23" />
                    <RANKING place="4" resultid="62" />
                    <RANKING place="1" resultid="169" />
                    <RANKING place="5" resultid="191" />
                    <RANKING place="6" resultid="202" />
                    <RANKING place="7" resultid="249" />
                    <RANKING place="2" resultid="414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="108" />
                    <RANKING place="6" resultid="164" />
                    <RANKING place="4" resultid="181" />
                    <RANKING place="3" resultid="392" />
                    <RANKING place="5" resultid="492" />
                    <RANKING place="7" resultid="503" />
                    <RANKING place="1" resultid="701" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="2" gender="M" round="PRE" order="2">
              <SWIMSTYLE name="100m Schmetterling männlich (Vorlauf)" stroke="FLY" relaycount="1" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="2001" number="1" daytime="10:08" />
                <HEAT heatid="2002" number="2" daytime="10:10" />
                <HEAT heatid="2003" number="3" daytime="10:12" />
                <HEAT heatid="2004" number="4" daytime="10:14" />
                <HEAT heatid="2005" number="5" daytime="10:16" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="306" />
                    <RANKING place="1" resultid="573" />
                    <RANKING place="3" resultid="667" />
                    <RANKING place="4" resultid="726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="96" />
                    <RANKING place="3" resultid="221" />
                    <RANKING place="6" resultid="590" />
                    <RANKING place="4" resultid="677" />
                    <RANKING place="5" resultid="721" />
                    <RANKING place="2" resultid="750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="8" resultid="12" />
                    <RANKING place="5" resultid="44" />
                    <RANKING place="1" resultid="102" />
                    <RANKING place="3" resultid="291" />
                    <RANKING place="4" resultid="553" />
                    <RANKING place="7" resultid="563" />
                    <RANKING place="2" resultid="579" />
                    <RANKING place="6" resultid="788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="144" />
                    <RANKING place="7" resultid="186" />
                    <RANKING place="1" resultid="364" />
                    <RANKING place="6" resultid="441" />
                    <RANKING place="5" resultid="455" />
                    <RANKING place="3" resultid="630" />
                    <RANKING place="8" resultid="682" />
                    <RANKING place="4" resultid="745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="134" />
                    <RANKING place="1" resultid="489" />
                    <RANKING place="4" resultid="737" />
                    <RANKING place="2" resultid="740" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="3" gender="F" round="TIM" order="3">
              <SWIMSTYLE name="200m Freistil weiblich" stroke="FREE" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="3001" number="1" daytime="10:18" />
                <HEAT heatid="3002" number="2" daytime="10:21" />
                <HEAT heatid="3003" number="3" daytime="10:24" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="315" />
                    <RANKING place="2" resultid="346" />
                    <RANKING place="3" resultid="778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="325" />
                    <RANKING place="2" resultid="340" />
                    <RANKING place="1" resultid="525" />
                    <RANKING place="3" resultid="774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="84" />
                    <RANKING place="3" resultid="208" />
                    <RANKING place="1" resultid="716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="281" />
                    <RANKING place="2" resultid="286" />
                    <RANKING place="1" resultid="520" />
                    <RANKING place="4" resultid="634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="73" />
                    <RANKING place="1" resultid="214" />
                    <RANKING place="3" resultid="218" />
                    <RANKING place="2" resultid="447" />
                    <RANKING place="5" resultid="513" />
                    <RANKING place="7" resultid="694" />
                    <RANKING place="6" resultid="702" />
                    <RANKING place="8" resultid="731" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="4" gender="M" round="TIM" order="4">
              <SWIMSTYLE name="200m Freistil männlich" stroke="FREE" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="4000" number="0" />
                <HEAT heatid="4001" number="1" daytime="10:27" />
                <HEAT heatid="4002" number="2" daytime="10:31" />
                <HEAT heatid="4003" number="3" daytime="10:34" />
                <HEAT heatid="4004" number="4" daytime="10:37" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="381" />
                    <RANKING place="2" resultid="485" />
                    <RANKING place="3" resultid="532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="227" />
                    <RANKING place="3" resultid="321" />
                    <RANKING place="4" resultid="496" />
                    <RANKING place="2" resultid="557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="78" />
                    <RANKING place="1" resultid="784" />
                    <RANKING place="3" resultid="798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="111" />
                    <RANKING place="4" resultid="296" />
                    <RANKING place="1" resultid="444" />
                    <RANKING place="3" resultid="481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="123" />
                    <RANKING place="3" resultid="244" />
                    <RANKING place="1" resultid="762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="9" resultid="8" />
                    <RANKING place="4" resultid="128" />
                    <RANKING place="2" resultid="242" />
                    <RANKING place="6" resultid="273" />
                    <RANKING place="1" resultid="278" />
                    <RANKING place="8" resultid="451" />
                    <RANKING place="7" resultid="467" />
                    <RANKING place="5" resultid="517" />
                    <RANKING place="3" resultid="734" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="5" gender="F" round="PRE" order="5">
              <SWIMSTYLE name="100m Brust weiblich (Vorlauf)" stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="5001" number="1" daytime="10:40" />
                <HEAT heatid="5002" number="2" daytime="10:43" />
                <HEAT heatid="5003" number="3" daytime="10:45" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="542" />
                    <RANKING place="2" resultid="756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="117" />
                    <RANKING place="2" resultid="547" />
                    <RANKING place="3" resultid="595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="5" resultid="24" />
                    <RANKING place="7" resultid="63" />
                    <RANKING place="4" resultid="90" />
                    <RANKING place="6" resultid="170" />
                    <RANKING place="3" resultid="387" />
                    <RANKING place="8" resultid="434" />
                    <RANKING place="1" resultid="463" />
                    <RANKING place="2" resultid="568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="35" />
                    <RANKING place="1" resultid="54" />
                    <RANKING place="3" resultid="352" />
                    <RANKING place="2" resultid="600" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="6" gender="M" round="PRE" order="6">
              <SWIMSTYLE name="100m Brust männlich (Vorlauf)" stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="6001" number="1" daytime="10:47" />
                <HEAT heatid="6002" number="2" daytime="10:50" />
                <HEAT heatid="6003" number="3" daytime="10:52" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="668" />
                    <RANKING place="1" resultid="727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="139" />
                    <RANKING place="3" resultid="232" />
                    <RANKING place="4" resultid="424" />
                    <RANKING place="6" resultid="591" />
                    <RANKING place="2" resultid="678" />
                    <RANKING place="5" resultid="722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="13" />
                    <RANKING place="1" resultid="310" />
                    <RANKING place="2" resultid="430" />
                    <RANKING place="3" resultid="564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="255" />
                    <RANKING place="2" resultid="473" />
                    <RANKING place="3" resultid="672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="68" />
                    <RANKING place="3" resultid="331" />
                    <RANKING place="1" resultid="355" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="7" gender="F" round="TIM" order="7">
              <SWIMSTYLE name="200m Rücken weiblich" stroke="BACK" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="7001" number="1" daytime="10:55" />
                <HEAT heatid="7002" number="2" daytime="10:59" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014" />
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="197" />
                    <RANKING place="2" resultid="341" />
                    <RANKING place="3" resultid="508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="335" />
                    <RANKING place="2" resultid="585" />
                    <RANKING place="1" resultid="626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="203" />
                    <RANKING place="6" resultid="250" />
                    <RANKING place="2" resultid="264" />
                    <RANKING place="4" resultid="287" />
                    <RANKING place="1" resultid="437" />
                    <RANKING place="5" resultid="659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="18" />
                    <RANKING place="1" resultid="165" />
                    <RANKING place="3" resultid="182" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="8" gender="M" round="TIM" order="8">
              <SWIMSTYLE name="200m Rücken männlich" stroke="BACK" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="8001" number="1" daytime="11:02" />
                <HEAT heatid="8002" number="2" daytime="11:06" />
                <HEAT heatid="8003" number="3" daytime="11:09" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="370" />
                    <RANKING place="2" resultid="486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="97" />
                    <RANKING place="3" resultid="425" />
                    <RANKING place="2" resultid="767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="79" />
                    <RANKING place="1" resultid="175" />
                    <RANKING place="3" resultid="800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="145" />
                    <RANKING place="2" resultid="187" />
                    <RANKING place="3" resultid="365" />
                    <RANKING place="4" resultid="664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="135" />
                    <RANKING place="1" resultid="401" />
                    <RANKING place="2" resultid="697" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="9" gender="F" round="TIM" order="9">
              <SWIMSTYLE name="800m Freistil weiblich" stroke="FREE" relaycount="1" distance="800" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="9000" number="0" />
                <HEAT heatid="9001" number="1" daytime="11:12" />
                <HEAT heatid="9002" number="2" daytime="11:24" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="689" />
                    <RANKING place="1" resultid="705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="613" />
                    <RANKING place="2" resultid="654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="209" />
                    <RANKING place="3" resultid="477" />
                    <RANKING place="2" resultid="608" />
                    <RANKING place="1" resultid="619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="219" />
                    <RANKING place="1" resultid="285" />
                    <RANKING place="3" resultid="695" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="10" number="10" gender="M" round="TIM" order="10">
              <SWIMSTYLE name="800m Freistil männlich" stroke="FREE" relaycount="1" distance="800" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="10000" number="0" />
                <HEAT heatid="10001" number="1" daytime="11:36" />
                <HEAT heatid="10002" number="2" daytime="11:48" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014" />
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="1" />
                    <RANKING place="2" resultid="29" />
                    <RANKING place="4" resultid="228" />
                    <RANKING place="1" resultid="359" />
                    <RANKING place="3" resultid="419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="5" resultid="39" />
                    <RANKING place="4" resultid="238" />
                    <RANKING place="3" resultid="376" />
                    <RANKING place="1" resultid="470" />
                    <RANKING place="2" resultid="785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011" />
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="57" />
                    <RANKING place="2" resultid="245" />
                    <RANKING place="4" resultid="631" />
                    <RANKING place="3" resultid="683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="5" />
                    <RANKING place="2" resultid="738" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="11" gender="F" round="PRE" order="11">
              <SWIMSTYLE name="100m Freistil weiblich (Vorlauf)" stroke="FREE" relaycount="1" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="11001" number="1" daytime="11:59" />
                <HEAT heatid="11002" number="2" daytime="12:01" />
                <HEAT heatid="11003" number="3" daytime="12:03" />
                <HEAT heatid="11004" number="4" daytime="12:04" />
                <HEAT heatid="11005" number="5" daytime="12:06" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="316" />
                    <RANKING place="2" resultid="347" />
                    <RANKING place="4" resultid="711" />
                    <RANKING place="3" resultid="779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="326" />
                    <RANKING place="2" resultid="526" />
                    <RANKING place="1" resultid="543" />
                    <RANKING place="3" resultid="757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="50" />
                    <RANKING place="3" resultid="85" />
                    <RANKING place="1" resultid="118" />
                    <RANKING place="5" resultid="548" />
                    <RANKING place="6" resultid="596" />
                    <RANKING place="4" resultid="717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="9" resultid="91" />
                    <RANKING place="6" resultid="171" />
                    <RANKING place="2" resultid="192" />
                    <RANKING place="11" resultid="268" />
                    <RANKING place="1" resultid="388" />
                    <RANKING place="4" resultid="405" />
                    <RANKING place="7" resultid="415" />
                    <RANKING place="3" resultid="438" />
                    <RANKING place="5" resultid="521" />
                    <RANKING place="8" resultid="569" />
                    <RANKING place="10" resultid="660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="74" />
                    <RANKING place="1" resultid="215" />
                    <RANKING place="2" resultid="260" />
                    <RANKING place="7" resultid="353" />
                    <RANKING place="4" resultid="393" />
                    <RANKING place="5" resultid="493" />
                    <RANKING place="6" resultid="504" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="12" number="12" gender="M" round="PRE" order="12">
              <SWIMSTYLE name="100m Freistil männlich (Vorlauf)" stroke="FREE" relaycount="1" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="12001" number="1" daytime="12:08" />
                <HEAT heatid="12002" number="2" daytime="12:10" />
                <HEAT heatid="12003" number="3" daytime="12:12" />
                <HEAT heatid="12004" number="4" daytime="12:13" />
                <HEAT heatid="12005" number="5" daytime="12:15" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="307" />
                    <RANKING place="2" resultid="371" />
                    <RANKING place="3" resultid="382" />
                    <RANKING place="5" resultid="533" />
                    <RANKING place="4" resultid="574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="222" />
                    <RANKING place="3" resultid="233" />
                    <RANKING place="7" resultid="322" />
                    <RANKING place="6" resultid="497" />
                    <RANKING place="4" resultid="558" />
                    <RANKING place="2" resultid="751" />
                    <RANKING place="5" resultid="768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="112" />
                    <RANKING place="4" resultid="292" />
                    <RANKING place="10" resultid="297" />
                    <RANKING place="5" resultid="311" />
                    <RANKING place="7" resultid="431" />
                    <RANKING place="1" resultid="445" />
                    <RANKING place="6" resultid="482" />
                    <RANKING place="9" resultid="539" />
                    <RANKING place="8" resultid="580" />
                    <RANKING place="3" resultid="789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="3" resultid="124" />
                    <RANKING place="4" resultid="256" />
                    <RANKING place="2" resultid="673" />
                    <RANKING place="5" resultid="746" />
                    <RANKING place="1" resultid="763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="10" resultid="9" />
                    <RANKING place="6" resultid="129" />
                    <RANKING place="7" resultid="274" />
                    <RANKING place="2" resultid="279" />
                    <RANKING place="8" resultid="452" />
                    <RANKING place="11" resultid="468" />
                    <RANKING place="1" resultid="490" />
                    <RANKING place="9" resultid="518" />
                    <RANKING place="5" resultid="698" />
                    <RANKING place="3" resultid="735" />
                    <RANKING place="4" resultid="741" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2025-07-05" daytime="01:30">
          <EVENTS>
            <EVENT eventid="13" number="101" gender="F" round="FIN" order="13">
              <SWIMSTYLE name="100m Schmetterling weiblich (Finale)" stroke="FLY" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="13001" number="1" daytime="13:47" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="15" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="803" />
                    <RANKING place="3" resultid="804" />
                    <RANKING place="4" resultid="805" />
                    <RANKING place="2" resultid="806" />
                    <RANKING place="6" resultid="807" />
                    <RANKING place="5" resultid="808" />
                    <RANKING place="7" resultid="809" />
                    <RANKING place="8" resultid="810" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="14" number="201" gender="F" round="FIN" order="14">
              <SWIMSTYLE name="100m Schmetterling weiblich (Finale)" stroke="FLY" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="14000" number="0" />
                <HEAT heatid="14001" number="1" daytime="13:49" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="16" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="813" />
                    <RANKING place="3" resultid="814" />
                    <RANKING place="5" resultid="815" />
                    <RANKING place="1" resultid="816" />
                    <RANKING place="4" resultid="817" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="15" number="102" gender="M" round="FIN" order="15">
              <SWIMSTYLE name="100m Schmetterling männlich (Finale)" stroke="FLY" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="15001" number="1" daytime="13:50" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="15" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="818" />
                    <RANKING place="1" resultid="819" />
                    <RANKING place="3" resultid="820" />
                    <RANKING place="4" resultid="821" />
                    <RANKING place="7" resultid="822" />
                    <RANKING place="8" resultid="823" />
                    <RANKING place="6" resultid="824" />
                    <RANKING place="5" resultid="825" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="16" number="202" gender="M" round="FIN" order="16">
              <SWIMSTYLE name="100m Schmetterling männlich (Finale)" stroke="FLY" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="16001" number="1" daytime="13:52" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="16" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="826" />
                    <RANKING place="2" resultid="827" />
                    <RANKING place="3" resultid="828" />
                    <RANKING place="4" resultid="829" />
                    <RANKING place="5" resultid="830" />
                    <RANKING place="6" resultid="831" />
                    <RANKING place="7" resultid="832" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="17" number="105" gender="F" round="FIN" order="17">
              <SWIMSTYLE name="100m Brust weiblich (Finale)" stroke="BREAST" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="17001" number="1" daytime="13:54" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="15" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="833" />
                    <RANKING place="4" resultid="834" />
                    <RANKING place="1" resultid="835" />
                    <RANKING place="3" resultid="836" />
                    <RANKING place="5" resultid="837" />
                    <RANKING place="7" resultid="838" />
                    <RANKING place="6" resultid="839" />
                    <RANKING place="8" resultid="840" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18" number="205" gender="F" round="FIN" order="18">
              <SWIMSTYLE name="100m Brust weiblich (Finale)" stroke="BREAST" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="18001" number="1" daytime="13:56" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="16" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="841" />
                    <RANKING place="2" resultid="842" />
                    <RANKING place="3" resultid="843" />
                    <RANKING place="4" resultid="844" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="19" number="106" gender="M" round="FIN" order="19">
              <SWIMSTYLE name="100m Brust männlich (Finale)" stroke="BREAST" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="19001" number="1" daytime="13:58" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="15" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="845" />
                    <RANKING place="3" resultid="846" />
                    <RANKING place="2" resultid="847" />
                    <RANKING place="4" resultid="848" />
                    <RANKING place="6" resultid="849" />
                    <RANKING place="5" resultid="850" />
                    <RANKING place="7" resultid="851" />
                    <RANKING place="8" resultid="852" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="20" number="206" gender="M" round="FIN" order="20">
              <SWIMSTYLE name="100m Brust männlich (Finale)" stroke="BREAST" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="20001" number="1" daytime="14:00" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="16" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="853" />
                    <RANKING place="2" resultid="854" />
                    <RANKING place="3" resultid="855" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="21" number="13" gender="F" round="TIM" order="21">
              <SWIMSTYLE name="50m Rücken weiblich" stroke="BACK" relaycount="1" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="21001" number="1" daytime="14:02" />
                <HEAT heatid="21002" number="2" daytime="14:03" />
                <HEAT heatid="21003" number="3" daytime="14:05" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="317" />
                    <RANKING place="1" resultid="348" />
                    <RANKING place="3" resultid="712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="342" />
                    <RANKING place="5" resultid="509" />
                    <RANKING place="3" resultid="527" />
                    <RANKING place="1" resultid="544" />
                    <RANKING place="4" resultid="758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="51" />
                    <RANKING place="2" resultid="210" />
                    <RANKING place="3" resultid="478" />
                    <RANKING place="4" resultid="549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="92" />
                    <RANKING place="2" resultid="265" />
                    <RANKING place="1" resultid="282" />
                    <RANKING place="5" resultid="288" />
                    <RANKING place="3" resultid="439" />
                    <RANKING place="6" resultid="522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="19" />
                    <RANKING place="3" resultid="36" />
                    <RANKING place="2" resultid="75" />
                    <RANKING place="1" resultid="220" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22" number="14" gender="M" round="TIM" order="22">
              <SWIMSTYLE name="50m Rücken männlich" stroke="BACK" relaycount="1" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="22001" number="1" daytime="14:06" />
                <HEAT heatid="22002" number="2" daytime="14:07" />
                <HEAT heatid="22003" number="3" daytime="14:08" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="372" />
                    <RANKING place="3" resultid="534" />
                    <RANKING place="2" resultid="575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="98" />
                    <RANKING place="5" resultid="140" />
                    <RANKING place="4" resultid="223" />
                    <RANKING place="2" resultid="234" />
                    <RANKING place="7" resultid="426" />
                    <RANKING place="6" resultid="559" />
                    <RANKING place="3" resultid="752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="239" />
                    <RANKING place="2" resultid="377" />
                    <RANKING place="1" resultid="412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="104" />
                    <RANKING place="2" resultid="483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="69" />
                    <RANKING place="2" resultid="130" />
                    <RANKING place="1" resultid="275" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23" number="15" gender="F" round="TIM" order="23">
              <SWIMSTYLE name="200m Lagen weiblich" stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="23001" number="1" daytime="14:10" />
                <HEAT heatid="23002" number="2" daytime="14:13" />
                <HEAT heatid="23003" number="3" daytime="14:17" />
                <HEAT heatid="23004" number="4" daytime="14:20" />
                <HEAT heatid="23005" number="5" daytime="14:24" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="3" resultid="318" />
                    <RANKING place="4" resultid="690" />
                    <RANKING place="2" resultid="706" />
                    <RANKING place="1" resultid="780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="198" />
                    <RANKING place="6" resultid="510" />
                    <RANKING place="4" resultid="528" />
                    <RANKING place="5" resultid="614" />
                    <RANKING place="3" resultid="655" />
                    <RANKING place="2" resultid="775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="7" resultid="86" />
                    <RANKING place="1" resultid="119" />
                    <RANKING place="5" resultid="154" />
                    <RANKING place="9" resultid="336" />
                    <RANKING place="2" resultid="397" />
                    <RANKING place="8" resultid="479" />
                    <RANKING place="3" resultid="586" />
                    <RANKING place="10" resultid="597" />
                    <RANKING place="4" resultid="620" />
                    <RANKING place="6" resultid="627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="25" />
                    <RANKING place="3" resultid="64" />
                    <RANKING place="5" resultid="193" />
                    <RANKING place="8" resultid="251" />
                    <RANKING place="6" resultid="269" />
                    <RANKING place="2" resultid="406" />
                    <RANKING place="4" resultid="416" />
                    <RANKING place="7" resultid="435" />
                    <RANKING place="10" resultid="635" />
                    <RANKING place="9" resultid="661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="55" />
                    <RANKING place="6" resultid="183" />
                    <RANKING place="3" resultid="261" />
                    <RANKING place="1" resultid="448" />
                    <RANKING place="4" resultid="514" />
                    <RANKING place="5" resultid="601" />
                    <RANKING place="7" resultid="732" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="24" number="16" gender="M" round="TIM" order="24">
              <SWIMSTYLE name="200m Lagen männlich" stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="24000" number="0" />
                <HEAT heatid="24001" number="1" daytime="14:27" />
                <HEAT heatid="24002" number="2" daytime="14:31" />
                <HEAT heatid="24003" number="3" daytime="14:34" />
                <HEAT heatid="24004" number="4" daytime="14:37" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="383" />
                    <RANKING place="3" resultid="487" />
                    <RANKING place="2" resultid="535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="7" resultid="2" />
                    <RANKING place="1" resultid="30" />
                    <RANKING place="4" resultid="323" />
                    <RANKING place="2" resultid="360" />
                    <RANKING place="3" resultid="420" />
                    <RANKING place="8" resultid="498" />
                    <RANKING place="6" resultid="560" />
                    <RANKING place="5" resultid="769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="40" />
                    <RANKING place="3" resultid="80" />
                    <RANKING place="2" resultid="177" />
                    <RANKING place="1" resultid="471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="14" />
                    <RANKING place="3" resultid="45" />
                    <RANKING place="1" resultid="113" />
                    <RANKING place="5" resultid="540" />
                    <RANKING place="2" resultid="554" />
                    <RANKING place="4" resultid="581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="58" />
                    <RANKING place="1" resultid="125" />
                    <RANKING place="4" resultid="188" />
                    <RANKING place="3" resultid="366" />
                    <RANKING place="5" resultid="684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="136" />
                    <RANKING place="1" resultid="243" />
                    <RANKING place="3" resultid="402" />
                    <RANKING place="2" resultid="699" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="25" number="17" gender="F" round="TIM" order="25">
              <SWIMSTYLE name="1500m Freistil weiblich" stroke="FREE" relaycount="1" distance="1500" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="25000" number="0" />
                <HEAT heatid="25001" number="1" daytime="14:40" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014" />
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="216" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26" number="18" gender="M" round="TIM" order="26">
              <SWIMSTYLE name="1500m Freistil männlich" stroke="FREE" relaycount="1" distance="1500" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="26001" number="1" daytime="15:01" />
                <HEAT heatid="26002" number="2" daytime="15:23" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="308" />
                    <RANKING place="2" resultid="669" />
                    <RANKING place="3" resultid="728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="229" />
                    <RANKING place="2" resultid="592" />
                    <RANKING place="4" resultid="679" />
                    <RANKING place="3" resultid="723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012" />
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="34" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="27" number="19" gender="F" round="TIM" order="27">
              <SWIMSTYLE name="50m Schmetterling weiblich" stroke="FLY" relaycount="1" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="27001" number="1" daytime="15:45" />
                <HEAT heatid="27002" number="2" daytime="15:47" />
                <HEAT heatid="27003" number="3" daytime="15:48" />
                <HEAT heatid="27004" number="4" daytime="15:49" />
                <HEAT heatid="27005" number="5" daytime="15:50" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="349" />
                    <RANKING place="2" resultid="713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="199" />
                    <RANKING place="4" resultid="343" />
                    <RANKING place="3" resultid="529" />
                    <RANKING place="2" resultid="545" />
                    <RANKING place="5" resultid="759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="87" />
                    <RANKING place="5" resultid="155" />
                    <RANKING place="6" resultid="211" />
                    <RANKING place="3" resultid="337" />
                    <RANKING place="2" resultid="398" />
                    <RANKING place="7" resultid="587" />
                    <RANKING place="8" resultid="609" />
                    <RANKING place="1" resultid="621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="26" />
                    <RANKING place="3" resultid="172" />
                    <RANKING place="7" resultid="252" />
                    <RANKING place="5" resultid="270" />
                    <RANKING place="1" resultid="389" />
                    <RANKING place="2" resultid="407" />
                    <RANKING place="6" resultid="464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="5" resultid="20" />
                    <RANKING place="1" resultid="56" />
                    <RANKING place="3" resultid="109" />
                    <RANKING place="4" resultid="166" />
                    <RANKING place="2" resultid="494" />
                    <RANKING place="6" resultid="505" />
                    <RANKING place="7" resultid="602" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="28" number="20" gender="M" round="TIM" order="28">
              <SWIMSTYLE name="50m Schmetterling männlich" stroke="FLY" relaycount="1" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="28001" number="1" daytime="15:51" />
                <HEAT heatid="28002" number="2" daytime="15:53" />
                <HEAT heatid="28003" number="3" daytime="15:54" />
                <HEAT heatid="28004" number="4" daytime="15:55" />
                <HEAT heatid="28005" number="5" daytime="15:57" />
                <HEAT heatid="28006" number="6" daytime="15:58" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="373" />
                    <RANKING place="3" resultid="488" />
                    <RANKING place="4" resultid="536" />
                    <RANKING place="1" resultid="576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="31" />
                    <RANKING place="3" resultid="224" />
                    <RANKING place="3" resultid="235" />
                    <RANKING place="8" resultid="324" />
                    <RANKING place="2" resultid="361" />
                    <RANKING place="7" resultid="421" />
                    <RANKING place="9" resultid="499" />
                    <RANKING place="1" resultid="753" />
                    <RANKING place="6" resultid="770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="5" resultid="41" />
                    <RANKING place="3" resultid="81" />
                    <RANKING place="2" resultid="178" />
                    <RANKING place="6" resultid="240" />
                    <RANKING place="4" resultid="378" />
                    <RANKING place="1" resultid="413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="15" />
                    <RANKING place="4" resultid="46" />
                    <RANKING place="1" resultid="114" />
                    <RANKING place="3" resultid="293" />
                    <RANKING place="5" resultid="298" />
                    <RANKING place="2" resultid="555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="7" resultid="59" />
                    <RANKING place="5" resultid="257" />
                    <RANKING place="1" resultid="367" />
                    <RANKING place="8" resultid="442" />
                    <RANKING place="4" resultid="456" />
                    <RANKING place="2" resultid="674" />
                    <RANKING place="9" resultid="685" />
                    <RANKING place="6" resultid="747" />
                    <RANKING place="2" resultid="764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="6" />
                    <RANKING place="6" resultid="10" />
                    <RANKING place="2" resultid="70" />
                    <RANKING place="5" resultid="491" />
                    <RANKING place="4" resultid="700" />
                    <RANKING place="7" resultid="739" />
                    <RANKING place="1" resultid="742" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="29" number="21" gender="F" round="TIM" order="29">
              <SWIMSTYLE name="200m Brust weiblich" stroke="BREAST" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="29001" number="1" daytime="15:59" />
                <HEAT heatid="29002" number="2" daytime="16:03" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="3" resultid="691" />
                    <RANKING place="2" resultid="707" />
                    <RANKING place="1" resultid="781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="615" />
                    <RANKING place="1" resultid="656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="120" />
                    <RANKING place="2" resultid="550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="65" />
                    <RANKING place="2" resultid="204" />
                    <RANKING place="4" resultid="436" />
                    <RANKING place="3" resultid="570" />
                    <RANKING place="5" resultid="636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="30" number="22" gender="M" round="TIM" order="30">
              <SWIMSTYLE name="200m Brust männlich" stroke="BREAST" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="30001" number="1" daytime="16:07" />
                <HEAT heatid="30002" number="2" daytime="16:11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="99" />
                    <RANKING place="2" resultid="141" />
                    <RANKING place="3" resultid="427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="105" />
                    <RANKING place="1" resultid="312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="146" />
                    <RANKING place="2" resultid="474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="131" />
                    <RANKING place="3" resultid="332" />
                    <RANKING place="1" resultid="356" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="31" number="111" gender="F" round="FIN" order="31">
              <SWIMSTYLE name="100m Freistil weiblich (Finale)" stroke="FREE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="31001" number="1" daytime="16:15" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="15" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="856" />
                    <RANKING place="3" resultid="857" />
                    <RANKING place="2" resultid="858" />
                    <RANKING place="5" resultid="859" />
                    <RANKING place="4" resultid="860" />
                    <RANKING place="6" resultid="861" />
                    <RANKING place="8" resultid="862" />
                    <RANKING place="7" resultid="863" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="32" number="211" gender="F" round="FIN" order="32">
              <SWIMSTYLE name="100m Freistil weiblich (Finale)" stroke="FREE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="32001" number="1" daytime="16:17" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="16" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="864" />
                    <RANKING place="2" resultid="865" />
                    <RANKING place="3" resultid="866" />
                    <RANKING place="4" resultid="867" />
                    <RANKING place="5" resultid="868" />
                    <RANKING place="6" resultid="869" />
                    <RANKING place="7" resultid="870" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="33" number="112" gender="M" round="FIN" order="33">
              <SWIMSTYLE name="100m Freistil männlich (Finale)" stroke="FREE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="33001" number="1" daytime="16:18" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="15" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="871" />
                    <RANKING place="2" resultid="872" />
                    <RANKING place="4" resultid="873" />
                    <RANKING place="3" resultid="874" />
                    <RANKING place="6" resultid="875" />
                    <RANKING place="5" resultid="876" />
                    <RANKING place="7" resultid="877" />
                    <RANKING place="8" resultid="878" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="34" number="212" gender="M" round="FIN" order="34">
              <SWIMSTYLE name="100m Freistil männlich (Finale)" stroke="FREE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="34000" number="0" />
                <HEAT heatid="34001" number="1" daytime="16:20" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="16" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="880" />
                    <RANKING place="2" resultid="881" />
                    <RANKING place="3" resultid="882" />
                    <RANKING place="4" resultid="883" />
                    <RANKING place="6" resultid="884" />
                    <RANKING place="8" resultid="885" />
                    <RANKING place="5" resultid="886" />
                    <RANKING place="7" resultid="887" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="3" date="2025-07-06" daytime="09:30" officialmeeting="09:00" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="35" number="23" gender="F" round="PRE" order="35">
              <SWIMSTYLE name="100m Rücken weiblich (Vorlauf)" stroke="BACK" relaycount="1" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="35001" number="1" daytime="09:30" />
                <HEAT heatid="35002" number="2" daytime="09:32" />
                <HEAT heatid="35003" number="3" daytime="09:34" />
                <HEAT heatid="35004" number="4" daytime="09:36" />
                <HEAT heatid="35005" number="5" daytime="09:38" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="692" />
                    <RANKING place="1" resultid="708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="200" />
                    <RANKING place="5" resultid="344" />
                    <RANKING place="7" resultid="511" />
                    <RANKING place="3" resultid="530" />
                    <RANKING place="4" resultid="616" />
                    <RANKING place="2" resultid="657" />
                    <RANKING place="6" resultid="760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="52" />
                    <RANKING place="3" resultid="121" />
                    <RANKING place="2" resultid="399" />
                    <RANKING place="6" resultid="598" />
                    <RANKING place="4" resultid="628" />
                    <RANKING place="5" resultid="719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="11" resultid="27" />
                    <RANKING place="5" resultid="94" />
                    <RANKING place="7" resultid="205" />
                    <RANKING place="13" resultid="253" />
                    <RANKING place="3" resultid="266" />
                    <RANKING place="12" resultid="271" />
                    <RANKING place="6" resultid="289" />
                    <RANKING place="1" resultid="390" />
                    <RANKING place="8" resultid="417" />
                    <RANKING place="2" resultid="440" />
                    <RANKING place="10" resultid="571" />
                    <RANKING place="14" resultid="637" />
                    <RANKING place="4" resultid="646" />
                    <RANKING place="9" resultid="662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="5" resultid="37" />
                    <RANKING place="2" resultid="76" />
                    <RANKING place="4" resultid="167" />
                    <RANKING place="1" resultid="262" />
                    <RANKING place="3" resultid="394" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="36" number="24" gender="M" round="PRE" order="36">
              <SWIMSTYLE name="100m Rücken männlich (Vorlauf)" stroke="BACK" relaycount="1" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="36001" number="1" daytime="09:40" />
                <HEAT heatid="36002" number="2" daytime="09:42" />
                <HEAT heatid="36003" number="3" daytime="09:44" />
                <HEAT heatid="36004" number="4" daytime="09:46" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="374" />
                    <RANKING place="4" resultid="537" />
                    <RANKING place="3" resultid="670" />
                    <RANKING place="2" resultid="729" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="100" />
                    <RANKING place="5" resultid="225" />
                    <RANKING place="7" resultid="428" />
                    <RANKING place="3" resultid="500" />
                    <RANKING place="4" resultid="593" />
                    <RANKING place="6" resultid="680" />
                    <RANKING place="2" resultid="724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="82" />
                    <RANKING place="2" resultid="801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="16" />
                    <RANKING place="5" resultid="47" />
                    <RANKING place="1" resultid="106" />
                    <RANKING place="4" resultid="115" />
                    <RANKING place="2" resultid="446" />
                    <RANKING place="3" resultid="541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="4" resultid="60" />
                    <RANKING place="2" resultid="247" />
                    <RANKING place="3" resultid="258" />
                    <RANKING place="5" resultid="368" />
                    <RANKING place="6" resultid="686" />
                    <RANKING place="1" resultid="765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="71" />
                    <RANKING place="5" resultid="137" />
                    <RANKING place="1" resultid="276" />
                    <RANKING place="4" resultid="357" />
                    <RANKING place="2" resultid="403" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="37" number="25" gender="F" round="TIM" order="37">
              <SWIMSTYLE name="200m Schmetterling weiblich" stroke="FLY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="37001" number="1" daytime="09:48" />
                <HEAT heatid="37002" number="2" daytime="09:52" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="350" />
                    <RANKING place="2" resultid="782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="156" />
                    <RANKING place="1" resultid="338" />
                    <RANKING place="3" resultid="588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="110" />
                    <RANKING place="2" resultid="184" />
                    <RANKING place="1" resultid="703" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="38" number="26" gender="M" round="TIM" order="38">
              <SWIMSTYLE name="200m Schmetterling männlich" stroke="FLY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="38001" number="1" daytime="09:56" />
                <HEAT heatid="38002" number="2" daytime="10:00" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014" />
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="294" />
                    <RANKING place="3" resultid="566" />
                    <RANKING place="2" resultid="582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="369" />
                    <RANKING place="3" resultid="443" />
                    <RANKING place="2" resultid="457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="7" />
                    <RANKING place="2" resultid="736" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="39" number="27" gender="F" round="TIM" order="39">
              <SWIMSTYLE name="50m Freistil weiblich" stroke="FREE" relaycount="1" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="39001" number="1" daytime="10:03" />
                <HEAT heatid="39002" number="2" daytime="10:05" />
                <HEAT heatid="39003" number="3" daytime="10:06" />
                <HEAT heatid="39004" number="4" daytime="10:07" />
                <HEAT heatid="39005" number="5" daytime="10:08" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="319" />
                    <RANKING place="3" resultid="714" />
                    <RANKING place="2" resultid="783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="53" />
                    <RANKING place="2" resultid="88" />
                    <RANKING place="6" resultid="212" />
                    <RANKING place="1" resultid="400" />
                    <RANKING place="7" resultid="551" />
                    <RANKING place="5" resultid="610" />
                    <RANKING place="3" resultid="622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="28" />
                    <RANKING place="6" resultid="173" />
                    <RANKING place="10" resultid="206" />
                    <RANKING place="9" resultid="272" />
                    <RANKING place="2" resultid="290" />
                    <RANKING place="4" resultid="391" />
                    <RANKING place="1" resultid="408" />
                    <RANKING place="7" resultid="418" />
                    <RANKING place="8" resultid="465" />
                    <RANKING place="5" resultid="523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="3" resultid="21" />
                    <RANKING place="6" resultid="77" />
                    <RANKING place="1" resultid="217" />
                    <RANKING place="4" resultid="263" />
                    <RANKING place="8" resultid="354" />
                    <RANKING place="7" resultid="395" />
                    <RANKING place="2" resultid="449" />
                    <RANKING place="5" resultid="495" />
                    <RANKING place="9" resultid="506" />
                    <RANKING place="10" resultid="515" />
                    <RANKING place="11" resultid="603" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="40" number="28" gender="M" round="TIM" order="40">
              <SWIMSTYLE name="50m Freistil männlich" stroke="FREE" relaycount="1" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="40000" number="0" />
                <HEAT heatid="40001" number="1" daytime="10:09" />
                <HEAT heatid="40002" number="2" daytime="10:10" />
                <HEAT heatid="40003" number="3" daytime="10:12" />
                <HEAT heatid="40004" number="4" daytime="10:13" />
                <HEAT heatid="40005" number="5" daytime="10:14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="375" />
                    <RANKING place="2" resultid="385" />
                    <RANKING place="3" resultid="577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="8" resultid="3" />
                    <RANKING place="4" resultid="32" />
                    <RANKING place="1" resultid="101" />
                    <RANKING place="7" resultid="142" />
                    <RANKING place="3" resultid="230" />
                    <RANKING place="9" resultid="422" />
                    <RANKING place="5" resultid="429" />
                    <RANKING place="2" resultid="754" />
                    <RANKING place="6" resultid="772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="42" />
                    <RANKING place="1" resultid="83" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="48" />
                    <RANKING place="2" resultid="107" />
                    <RANKING place="5" resultid="299" />
                    <RANKING place="3" resultid="313" />
                    <RANKING place="1" resultid="432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="8" resultid="61" />
                    <RANKING place="3" resultid="126" />
                    <RANKING place="1" resultid="147" />
                    <RANKING place="5" resultid="189" />
                    <RANKING place="6" resultid="632" />
                    <RANKING place="4" resultid="675" />
                    <RANKING place="7" resultid="748" />
                    <RANKING place="2" resultid="766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="7" resultid="11" />
                    <RANKING place="3" resultid="132" />
                    <RANKING place="6" resultid="138" />
                    <RANKING place="4" resultid="277" />
                    <RANKING place="1" resultid="454" />
                    <RANKING place="5" resultid="469" />
                    <RANKING place="2" resultid="743" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="41" number="29" gender="F" round="TIM" order="41">
              <SWIMSTYLE name="400m Lagen weiblich" stroke="MEDLEY" relaycount="1" distance="400" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="41000" number="0" />
                <HEAT heatid="41001" number="1" daytime="10:15" />
                <HEAT heatid="41002" number="2" daytime="10:23" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="3" resultid="351" />
                    <RANKING place="2" resultid="693" />
                    <RANKING place="1" resultid="709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="201" />
                    <RANKING place="4" resultid="345" />
                    <RANKING place="3" resultid="617" />
                    <RANKING place="2" resultid="658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="480" />
                    <RANKING place="2" resultid="629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="66" />
                    <RANKING place="3" resultid="638" />
                    <RANKING place="1" resultid="647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="696" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="42" number="30" gender="M" round="TIM" order="42">
              <SWIMSTYLE name="400m Lagen männlich" stroke="MEDLEY" relaycount="1" distance="400" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="42000" number="0" />
                <HEAT heatid="42001" number="1" daytime="10:30" />
                <HEAT heatid="42002" number="2" daytime="10:37" />
                <HEAT heatid="42003" number="3" daytime="10:44" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="309" />
                    <RANKING place="2" resultid="386" />
                    <RANKING place="3" resultid="671" />
                    <RANKING place="4" resultid="730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="226" />
                    <RANKING place="3" resultid="231" />
                    <RANKING place="5" resultid="594" />
                    <RANKING place="2" resultid="681" />
                    <RANKING place="4" resultid="725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="116" />
                    <RANKING place="3" resultid="484" />
                    <RANKING place="2" resultid="556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="475" />
                    <RANKING place="1" resultid="666" />
                    <RANKING place="3" resultid="687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="43" number="31" gender="F" round="TIM" order="43">
              <SWIMSTYLE name="50m Brust weiblich" stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="43001" number="1" daytime="10:51" />
                <HEAT heatid="43002" number="2" daytime="10:52" />
                <HEAT heatid="43003" number="3" daytime="10:54" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="122" />
                    <RANKING place="2" resultid="157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="95" />
                    <RANKING place="4" resultid="207" />
                    <RANKING place="2" resultid="284" />
                    <RANKING place="6" resultid="466" />
                    <RANKING place="5" resultid="524" />
                    <RANKING place="1" resultid="572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter">
                  <RANKINGS>
                    <RANKING place="5" resultid="22" />
                    <RANKING place="3" resultid="38" />
                    <RANKING place="4" resultid="168" />
                    <RANKING place="6" resultid="185" />
                    <RANKING place="1" resultid="450" />
                    <RANKING place="7" resultid="516" />
                    <RANKING place="2" resultid="604" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="44" number="32" gender="M" round="TIM" order="44">
              <SWIMSTYLE name="50m Brust männlich" stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="44000" number="0" />
                <HEAT heatid="44001" number="1" daytime="10:55" />
                <HEAT heatid="44002" number="2" daytime="10:56" />
                <HEAT heatid="44003" number="3" daytime="10:58" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="237" />
                    <RANKING place="3" resultid="501" />
                    <RANKING place="1" resultid="755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="17" />
                    <RANKING place="1" resultid="433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="259" />
                    <RANKING place="4" resultid="458" />
                    <RANKING place="2" resultid="633" />
                    <RANKING place="3" resultid="749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="72" />
                    <RANKING place="6" resultid="133" />
                    <RANKING place="3" resultid="333" />
                    <RANKING place="1" resultid="358" />
                    <RANKING place="5" resultid="404" />
                    <RANKING place="4" resultid="744" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="45" number="33" gender="F" round="TIM" order="45">
              <SWIMSTYLE name="400m Freistil weiblich" stroke="FREE" relaycount="1" distance="400" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="45001" number="1" daytime="10:59" />
                <HEAT heatid="45002" number="2" daytime="11:06" />
                <HEAT heatid="45003" number="3" daytime="11:12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="512" />
                    <RANKING place="1" resultid="531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="6" resultid="89" />
                    <RANKING place="7" resultid="213" />
                    <RANKING place="5" resultid="339" />
                    <RANKING place="8" resultid="552" />
                    <RANKING place="4" resultid="589" />
                    <RANKING place="9" resultid="599" />
                    <RANKING place="3" resultid="611" />
                    <RANKING place="2" resultid="623" />
                    <RANKING place="1" resultid="720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="67" />
                    <RANKING place="1" resultid="174" />
                    <RANKING place="5" resultid="254" />
                    <RANKING place="2" resultid="409" />
                    <RANKING place="4" resultid="663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="16" name="Jahrgang 2009 und älter" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="46" number="34" gender="M" round="TIM" order="46">
              <SWIMSTYLE name="400m Freistil männlich" stroke="FREE" relaycount="1" distance="400" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="46000" number="0" />
                <HEAT heatid="46001" number="1" daytime="11:18" />
                <HEAT heatid="46002" number="2" daytime="11:25" />
                <HEAT heatid="46003" number="3" daytime="11:30" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="11" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="12" agemin="12" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="4" />
                    <RANKING place="1" resultid="33" />
                    <RANKING place="2" resultid="143" />
                    <RANKING place="3" resultid="423" />
                    <RANKING place="5" resultid="502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="13" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="43" />
                    <RANKING place="2" resultid="241" />
                    <RANKING place="1" resultid="787" />
                    <RANKING place="4" resultid="802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="14" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="300" />
                    <RANKING place="3" resultid="314" />
                    <RANKING place="4" resultid="567" />
                    <RANKING place="1" resultid="583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="16" agemin="15" name="Jahrgang 2009/2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="127" />
                    <RANKING place="1" resultid="148" />
                    <RANKING place="4" resultid="190" />
                    <RANKING place="3" resultid="248" />
                    <RANKING place="5" resultid="676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="17" name="Jahrgang 2008 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="280" />
                    <RANKING place="2" resultid="519" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="47" number="123" gender="F" round="FIN" order="47">
              <SWIMSTYLE name="100m Rücken weiblich (Finale)" stroke="BACK" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="47001" number="1" daytime="11:36" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="15" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="888" />
                    <RANKING place="4" resultid="889" />
                    <RANKING place="3" resultid="890" />
                    <RANKING place="7" resultid="891" />
                    <RANKING place="5" resultid="892" />
                    <RANKING place="2" resultid="893" />
                    <RANKING place="6" resultid="894" />
                    <RANKING place="8" resultid="895" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="48" number="223" gender="F" round="FIN" order="48">
              <SWIMSTYLE name="100m Rücken weiblich (Finale)" stroke="BACK" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="48001" number="1" daytime="11:38" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="16" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="896" />
                    <RANKING place="2" resultid="897" />
                    <RANKING place="4" resultid="898" />
                    <RANKING place="3" resultid="899" />
                    <RANKING place="5" resultid="900" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="49" number="124" gender="M" round="FIN" order="49">
              <SWIMSTYLE name="100m Rücken männlich (Finale)" stroke="BACK" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="49001" number="1" daytime="11:40" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="15" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="901" />
                    <RANKING place="2" resultid="902" />
                    <RANKING place="4" resultid="903" />
                    <RANKING place="3" resultid="904" />
                    <RANKING place="5" resultid="905" />
                    <RANKING place="7" resultid="906" />
                    <RANKING place="6" resultid="907" />
                    <RANKING place="8" resultid="908" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="50" number="224" gender="M" round="FIN" order="50">
              <SWIMSTYLE name="100m Rücken männlich (Finale)" stroke="BACK" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="50001" number="1" daytime="11:41" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="16" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="909" />
                    <RANKING place="3" resultid="910" />
                    <RANKING place="2" resultid="911" />
                    <RANKING place="7" resultid="912" />
                    <RANKING place="8" resultid="913" />
                    <RANKING place="4" resultid="914" />
                    <RANKING place="5" resultid="915" />
                    <RANKING place="6" resultid="916" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="ATSV Freiberg e.V." nation="GER" region="12" code="3324">
          <ATHLETES>
            <ATHLETE athleteid="65" birthdate="2011-01-01" gender="M" lastname="Rehman" firstname="Roshan" license="431996" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:13.56" heatid="6001" lane="5" />
                <ENTRY eventid="12" entrytime="00:01:00.01" heatid="12005" lane="8" />
                <ENTRY eventid="30" entrytime="00:02:40.06" heatid="30002" lane="7" />
                <ENTRY eventid="40" entrytime="00:00:27.46" heatid="40004" lane="8" />
                <ENTRY eventid="46" entrytime="00:04:44.28" heatid="46002" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:14.34" heatid="19001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="310" eventid="6" swimtime="00:01:14.34" lane="5" heatid="6001" points="447" />
                <RESULT resultid="311" eventid="12" swimtime="00:00:59.84" lane="8" heatid="12005" points="466" />
                <RESULT resultid="847" eventid="19" swimtime="00:01:12.70" lane="3" heatid="19001" points="478" />
                <RESULT resultid="312" eventid="30" swimtime="00:02:43.31" lane="7" heatid="30002" points="453">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="313" eventid="40" swimtime="00:00:28.10" lane="8" heatid="40004" points="412" />
                <RESULT resultid="314" eventid="46" swimtime="00:04:45.82" lane="4" heatid="46002" points="456">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.48" />
                    <SPLIT distance="200" swimtime="00:02:19.77" />
                    <SPLIT distance="300" swimtime="00:03:33.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="DLRG Ortsgruppe Wernigerode" nation="GER" region="13" code="7154">
          <ATHLETES>
            <ATHLETE athleteid="156" birthdate="2009-01-01" gender="F" lastname="Vasic" firstname="Magdalena" license="396823" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:19.93" heatid="3002" lane="2" />
                <ENTRY eventid="23" entrytime="00:02:36.31" heatid="23004" lane="7" />
                <ENTRY eventid="45" entrytime="00:04:48.88" heatid="45003" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="731" eventid="3" swimtime="00:02:22.41" lane="2" heatid="3002" points="489">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="732" eventid="23" swimtime="00:02:42.94" lane="7" heatid="23004" points="463">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="733" eventid="45" status="WDR" swimtime="00:00:00.00" lane="5" heatid="45003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Dresdner Delphine e.V." nation="GER" region="12" code="5753">
          <ATHLETES>
            <ATHLETE athleteid="162" birthdate="2013-01-01" gender="F" lastname="Böhmert" firstname="Charlotte Katrin" license="437495" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:39.61" heatid="5003" lane="7" />
                <ENTRY eventid="11" entrytime="00:01:15.03" heatid="11001" lane="5" />
                <ENTRY eventid="21" entrytime="00:00:39.70" heatid="21001" lane="5" />
                <ENTRY eventid="27" entrytime="00:00:38.00" heatid="27002" lane="7" />
                <ENTRY eventid="35" entrytime="00:01:25.56" heatid="35002" lane="8" />
                <ENTRY eventid="39" entrytime="00:00:34.32" heatid="39001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="756" eventid="5" swimtime="00:01:37.16" lane="7" heatid="5003" points="287" />
                <RESULT resultid="757" eventid="11" swimtime="00:01:13.86" lane="5" heatid="11001" points="343" />
                <RESULT resultid="758" eventid="21" swimtime="00:00:38.46" lane="5" heatid="21001" points="340" />
                <RESULT resultid="759" eventid="27" swimtime="00:00:37.15" lane="7" heatid="27002" points="284" />
                <RESULT resultid="760" eventid="35" swimtime="00:01:25.51" lane="8" heatid="35002" points="298" />
                <RESULT resultid="761" eventid="39" swimtime="00:00:33.83" lane="5" heatid="39001" points="339" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163" birthdate="2009-01-01" gender="M" lastname="Müller" firstname="Emil" license="395288" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:00.09" heatid="4004" lane="2" />
                <ENTRY eventid="12" entrytime="00:00:55.52" heatid="12003" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:27.90" heatid="28005" lane="5" />
                <ENTRY eventid="36" entrytime="00:01:03.92" heatid="36002" lane="5" />
                <ENTRY eventid="40" entrytime="00:00:25.44" heatid="40005" lane="7" />
                <ENTRY eventid="50" entrytime="00:01:05.68" heatid="50001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="762" eventid="4" swimtime="00:02:03.09" lane="2" heatid="4004" points="569">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="763" eventid="12" swimtime="00:00:57.06" lane="3" heatid="12003" points="537" />
                <RESULT resultid="764" eventid="28" swimtime="00:00:28.15" lane="5" heatid="28005" points="495" />
                <RESULT resultid="765" eventid="36" swimtime="00:01:05.68" lane="5" heatid="36002" points="484" />
                <RESULT resultid="766" eventid="40" swimtime="00:00:26.61" lane="7" heatid="40005" points="485" />
                <RESULT resultid="912" eventid="50" swimtime="00:01:05.91" lane="6" heatid="50001" points="479" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164" birthdate="2013-01-01" gender="M" lastname="Böhmert" firstname="Flinn Jan" license="437496" nation="GER">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:02:52.32" heatid="8001" lane="4" />
                <ENTRY eventid="12" entrytime="00:01:12.16" heatid="12001" lane="3" />
                <ENTRY eventid="24" entrytime="00:02:56.09" heatid="24001" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:35.41" heatid="28002" lane="6" />
                <ENTRY eventid="38" entrytime="00:03:35.34" heatid="38001" lane="2" />
                <ENTRY eventid="40" entrytime="00:00:32.96" heatid="40001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="767" eventid="8" swimtime="00:02:49.97" lane="4" heatid="8001" points="285">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="768" eventid="12" swimtime="00:01:10.36" lane="3" heatid="12001" points="286" />
                <RESULT resultid="769" eventid="24" swimtime="00:02:55.45" lane="3" heatid="24001" points="274">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="770" eventid="28" swimtime="00:00:35.23" lane="6" heatid="28002" points="252" />
                <RESULT resultid="771" eventid="38" swimtime="00:03:14.34" lane="2" heatid="38001" points="183">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="772" eventid="40" swimtime="00:00:31.93" lane="6" heatid="40001" points="280" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165" birthdate="2013-01-01" gender="F" lastname="Hänig" firstname="Jasna" license="445403" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:14.49" heatid="1003" lane="8" />
                <ENTRY eventid="3" entrytime="00:02:30.14" heatid="3002" lane="8" />
                <ENTRY eventid="23" entrytime="00:02:45.24" heatid="23002" lane="3" />
                <ENTRY eventid="37" entrytime="00:02:50.77" heatid="37002" lane="2" />
                <ENTRY eventid="43" entrytime="00:00:41.36" heatid="43002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="773" eventid="1" swimtime="00:01:15.70" lane="8" heatid="1003" points="387" />
                <RESULT resultid="774" eventid="3" swimtime="00:02:35.99" lane="8" heatid="3002" points="372">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="775" eventid="23" swimtime="00:02:46.33" lane="3" heatid="23002" points="435">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="776" eventid="37" swimtime="00:03:03.12" lane="2" heatid="37002" points="294">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="777" eventid="43" swimtime="00:00:43.50" lane="1" heatid="43002" points="301" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166" birthdate="2014-01-01" gender="F" lastname="Richter" firstname="Marie-Sophie" license="447792" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:46.92" heatid="3001" lane="1" />
                <ENTRY eventid="11" entrytime="00:01:14.57" heatid="11002" lane="7" />
                <ENTRY eventid="23" entrytime="00:02:51.22" heatid="23002" lane="8" />
                <ENTRY eventid="29" entrytime="00:03:11.51" heatid="29002" lane="1" />
                <ENTRY eventid="37" entrytime="00:03:25.37" heatid="37001" lane="3" />
                <ENTRY eventid="39" entrytime="00:00:33.11" heatid="39002" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="778" eventid="3" swimtime="00:02:40.01" lane="1" heatid="3001" points="345">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="779" eventid="11" swimtime="00:01:13.89" lane="7" heatid="11002" points="342" />
                <RESULT resultid="780" eventid="23" swimtime="00:02:49.66" lane="8" heatid="23002" points="410">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="781" eventid="29" swimtime="00:03:08.18" lane="1" heatid="29002" points="390">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="782" eventid="37" swimtime="00:03:15.40" lane="3" heatid="37001" points="242">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="783" eventid="39" swimtime="00:00:33.23" lane="8" heatid="39002" points="358" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="2012-01-01" gender="M" lastname="Haberkorn" firstname="Matthäus" license="437400" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:15.79" heatid="4002" lane="4" />
                <ENTRY eventid="10" entrytime="00:09:27.51" heatid="10002" lane="2" />
                <ENTRY eventid="30" entrytime="00:02:46.89" heatid="30002" lane="8" />
                <ENTRY eventid="46" entrytime="00:04:46.16" heatid="46002" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="784" eventid="4" swimtime="00:02:14.71" lane="4" heatid="4002" points="434">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="785" eventid="10" swimtime="00:09:40.54" lane="2" heatid="10002" points="472">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="200" swimtime="00:02:17.97" />
                    <SPLIT distance="300" swimtime="00:03:30.37" />
                    <SPLIT distance="400" swimtime="00:04:44.47" />
                    <SPLIT distance="500" swimtime="00:05:59.38" />
                    <SPLIT distance="600" swimtime="00:07:13.43" />
                    <SPLIT distance="700" swimtime="00:08:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="786" eventid="30" swimtime="00:02:52.92" lane="8" heatid="30002" points="382">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="787" eventid="46" swimtime="00:04:41.07" lane="5" heatid="46002" points="479">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="200" swimtime="00:02:16.72" />
                    <SPLIT distance="300" swimtime="00:03:29.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="168" birthdate="2011-01-01" gender="M" lastname="Gennerich" firstname="Maximilian" license="423096" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:04.45" heatid="2003" lane="6" />
                <ENTRY eventid="12" entrytime="00:00:58.82" heatid="12004" lane="7" />
                <ENTRY eventid="38" entrytime="00:03:01.81" heatid="38001" lane="6" />
                <ENTRY eventid="42" entrytime="00:05:33.46" heatid="42000" lane="0" />
                <ENTRY eventid="33" entrytime="00:00:59.34" heatid="33001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="788" eventid="2" swimtime="00:01:07.48" lane="6" heatid="2003" points="393" />
                <RESULT resultid="789" eventid="12" swimtime="00:00:59.34" lane="7" heatid="12004" points="478" />
                <RESULT resultid="876" eventid="33" swimtime="00:00:58.88" lane="7" heatid="33001" points="489" />
                <RESULT resultid="790" eventid="38" status="WDR" swimtime="00:00:00.00" lane="6" heatid="38001" />
                <RESULT resultid="791" eventid="42" status="WDR" swimtime="00:00:00.00" lane="0" heatid="42000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169" birthdate="2012-01-01" gender="F" lastname="Müller" firstname="Milene" license="437414" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:23.83" heatid="5001" lane="6" />
                <ENTRY eventid="23" entrytime="00:02:45.69" heatid="23002" lane="6" />
                <ENTRY eventid="29" entrytime="00:03:02.69" heatid="29002" lane="7" />
                <ENTRY eventid="35" entrytime="00:01:16.12" heatid="35003" lane="8" />
                <ENTRY eventid="39" entrytime="00:00:29.80" heatid="39002" lane="5" />
                <ENTRY eventid="43" entrytime="00:00:37.53" heatid="43003" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="792" eventid="5" status="DNS" swimtime="00:00:00.00" lane="6" heatid="5001" />
                <RESULT resultid="793" eventid="23" status="DNS" swimtime="00:00:00.00" lane="6" heatid="23002" />
                <RESULT resultid="794" eventid="29" status="DNS" swimtime="00:00:00.00" lane="7" heatid="29002" />
                <RESULT resultid="795" eventid="35" status="DNS" swimtime="00:00:00.00" lane="8" heatid="35003" />
                <RESULT resultid="796" eventid="39" status="DNS" swimtime="00:00:00.00" lane="5" heatid="39002" />
                <RESULT resultid="797" eventid="43" status="DNS" swimtime="00:00:00.00" lane="8" heatid="43003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Dresdner SC 1898" nation="GER" region="12" code="3332">
          <ATHLETES>
            <ATHLETE athleteid="69" birthdate="2008-01-01" gender="M" lastname="Zische" firstname="Adrian" license="380817" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:05.39" heatid="6001" lane="4" />
                <ENTRY eventid="30" entrytime="00:02:22.54" heatid="30002" lane="5" />
                <ENTRY eventid="44" entrytime="00:00:30.21" heatid="44003" lane="5" />
                <ENTRY eventid="20" entrytime="00:01:10.97" heatid="20001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="331" eventid="6" swimtime="00:01:10.97" lane="4" heatid="6001" points="514" />
                <RESULT resultid="855" eventid="20" swimtime="00:01:10.30" lane="3" heatid="20001" points="529" />
                <RESULT resultid="332" eventid="30" swimtime="00:02:40.21" lane="5" heatid="30002" points="480">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="333" eventid="44" swimtime="00:00:31.95" lane="5" heatid="44003" points="535" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="70" birthdate="2012-01-01" gender="F" lastname="Kirberger" firstname="Alexandra" license="436906" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:11.65" heatid="1003" lane="7" />
                <ENTRY eventid="7" entrytime="00:02:39.81" heatid="7001" lane="4" />
                <ENTRY eventid="23" entrytime="00:02:44.14" heatid="23003" lane="8" />
                <ENTRY eventid="27" entrytime="00:00:30.92" heatid="27004" lane="6" />
                <ENTRY eventid="37" entrytime="00:02:40.82" heatid="37002" lane="6" />
                <ENTRY eventid="45" entrytime="00:05:09.00" heatid="45003" lane="8" />
                <ENTRY eventid="13" entrytime="00:01:10.64" heatid="13001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="334" eventid="1" swimtime="00:01:10.64" lane="7" heatid="1003" points="476" />
                <RESULT resultid="335" eventid="7" swimtime="00:02:39.87" lane="4" heatid="7001" points="456">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="807" eventid="13" swimtime="00:01:10.90" lane="2" heatid="13001" points="471" />
                <RESULT resultid="336" eventid="23" swimtime="00:02:43.26" lane="8" heatid="23003" points="461">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="337" eventid="27" swimtime="00:00:31.54" lane="6" heatid="27004" points="464" />
                <RESULT resultid="338" eventid="37" swimtime="00:02:44.67" lane="6" heatid="37002" points="404">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="339" eventid="45" swimtime="00:05:08.53" lane="8" heatid="45003" points="444">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.73" />
                    <SPLIT distance="200" swimtime="00:02:31.34" />
                    <SPLIT distance="300" swimtime="00:03:51.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="71" birthdate="2013-01-01" gender="F" lastname="Schwendler" firstname="Alexandra" license="449958" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:39.57" heatid="3001" lane="3" />
                <ENTRY eventid="7" entrytime="00:02:54.67" heatid="7001" lane="6" />
                <ENTRY eventid="21" entrytime="00:00:38.00" heatid="21001" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:35.30" heatid="27002" lane="6" />
                <ENTRY eventid="35" entrytime="00:01:19.41" heatid="35002" lane="6" />
                <ENTRY eventid="41" entrytime="00:06:40.44" heatid="41002" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="340" eventid="3" swimtime="00:02:35.40" lane="3" heatid="3001" points="376">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="341" eventid="7" swimtime="00:02:54.81" lane="6" heatid="7001" points="349">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="342" eventid="21" swimtime="00:00:37.05" lane="4" heatid="21001" points="381" />
                <RESULT resultid="343" eventid="27" swimtime="00:00:36.53" lane="6" heatid="27002" points="299" />
                <RESULT resultid="344" eventid="35" swimtime="00:01:23.54" lane="6" heatid="35002" points="319" />
                <RESULT resultid="345" eventid="41" swimtime="00:06:20.66" lane="8" heatid="41002" points="335">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.76" />
                    <SPLIT distance="200" swimtime="00:03:03.08" />
                    <SPLIT distance="300" swimtime="00:04:56.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="72" birthdate="2014-01-01" gender="F" lastname="Gutjahr" firstname="Anna Lena" license="448021" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:39.61" heatid="3001" lane="6" />
                <ENTRY eventid="11" entrytime="00:01:12.99" heatid="11002" lane="6" />
                <ENTRY eventid="21" entrytime="00:00:35.99" heatid="21002" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:33.99" heatid="27002" lane="4" />
                <ENTRY eventid="37" entrytime="00:02:57.21" heatid="37002" lane="8" />
                <ENTRY eventid="41" entrytime="00:06:50.92" heatid="41001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="346" eventid="3" swimtime="00:02:39.65" lane="6" heatid="3001" points="347">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="347" eventid="11" swimtime="00:01:13.39" lane="6" heatid="11002" points="349" />
                <RESULT resultid="348" eventid="21" swimtime="00:00:36.41" lane="2" heatid="21002" points="401" />
                <RESULT resultid="349" eventid="27" swimtime="00:00:33.01" lane="4" heatid="27002" points="405" />
                <RESULT resultid="350" eventid="37" swimtime="00:03:01.05" lane="8" heatid="37002" points="304">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="351" eventid="41" swimtime="00:06:23.20" lane="4" heatid="41001" points="328">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.48" />
                    <SPLIT distance="200" swimtime="00:03:01.62" />
                    <SPLIT distance="300" swimtime="00:04:56.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="73" birthdate="2009-01-01" gender="F" lastname="Zische" firstname="Annika" license="393879" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:12.93" heatid="5001" lane="4" />
                <ENTRY eventid="11" entrytime="00:01:00.59" heatid="11005" lane="3" />
                <ENTRY eventid="39" entrytime="00:00:27.39" heatid="39005" lane="1" />
                <ENTRY eventid="18" entrytime="00:01:16.14" heatid="18001" lane="3" />
                <ENTRY eventid="32" entrytime="00:01:02.97" heatid="32001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="352" eventid="5" swimtime="00:01:16.14" lane="4" heatid="5001" points="597" />
                <RESULT resultid="353" eventid="11" swimtime="00:01:02.97" lane="3" heatid="11005" points="553" />
                <RESULT resultid="843" eventid="18" swimtime="00:01:16.01" lane="3" heatid="18001" points="600" />
                <RESULT resultid="870" eventid="32" swimtime="00:01:03.33" lane="1" heatid="32001" points="544" />
                <RESULT resultid="354" eventid="39" swimtime="00:00:28.65" lane="1" heatid="39005" points="559" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="74" birthdate="2006-01-01" gender="M" lastname="Wüstenhagen" firstname="Arian" license="349848" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:01.05" heatid="6003" lane="4" />
                <ENTRY eventid="30" entrytime="00:02:16.91" heatid="30002" lane="4" />
                <ENTRY eventid="36" entrytime="00:01:04.29" heatid="36004" lane="3" />
                <ENTRY eventid="44" entrytime="00:00:28.06" heatid="44003" lane="4" />
                <ENTRY eventid="20" entrytime="00:01:02.82" heatid="20001" lane="4" />
                <ENTRY eventid="50" entrytime="00:01:06.73" heatid="50001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="355" eventid="6" swimtime="00:01:02.82" lane="4" heatid="6003" points="742" />
                <RESULT resultid="853" eventid="20" swimtime="00:01:03.06" lane="4" heatid="20001" points="733" />
                <RESULT resultid="356" eventid="30" swimtime="00:02:25.65" lane="4" heatid="30002" points="639">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="357" eventid="36" swimtime="00:01:06.73" lane="3" heatid="36004" points="462" />
                <RESULT resultid="358" eventid="44" swimtime="00:00:28.80" lane="4" heatid="44003" points="731" />
                <RESULT resultid="914" eventid="50" swimtime="00:01:02.83" lane="7" heatid="50001" points="553" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="75" birthdate="2013-01-01" gender="M" lastname="Lange" firstname="Arthur" license="443672" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:10:38.60" heatid="10001" lane="3" />
                <ENTRY eventid="24" entrytime="00:02:42.24" heatid="24002" lane="7" />
                <ENTRY eventid="28" entrytime="00:00:33.22" heatid="28003" lane="7" />
                <ENTRY eventid="40" entrytime="00:00:30.89" heatid="40002" lane="2" />
                <ENTRY eventid="46" entrytime="00:05:01.88" heatid="46000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="359" eventid="10" swimtime="00:10:28.92" lane="3" heatid="10001" points="371">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="200" swimtime="00:02:30.37" />
                    <SPLIT distance="300" swimtime="00:03:50.39" />
                    <SPLIT distance="400" swimtime="00:05:11.44" />
                    <SPLIT distance="500" swimtime="00:06:32.25" />
                    <SPLIT distance="600" swimtime="00:07:52.72" />
                    <SPLIT distance="700" swimtime="00:09:12.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="360" eventid="24" swimtime="00:02:42.18" lane="7" heatid="24002" points="347">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="361" eventid="28" swimtime="00:00:32.95" lane="7" heatid="28003" points="308" />
                <RESULT resultid="362" eventid="40" status="WDR" swimtime="00:00:00.00" lane="2" heatid="40002" />
                <RESULT resultid="363" eventid="46" status="WDR" swimtime="00:00:00.00" lane="0" heatid="46000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="76" birthdate="2009-01-01" gender="M" lastname="Wüstenhagen" firstname="Aurel" license="395576" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:00:59.37" heatid="2004" lane="5" />
                <ENTRY eventid="8" entrytime="00:02:28.31" heatid="8002" lane="3" />
                <ENTRY eventid="24" entrytime="00:02:22.51" heatid="24004" lane="8" />
                <ENTRY eventid="28" entrytime="00:00:27.10" heatid="28006" lane="7" />
                <ENTRY eventid="36" entrytime="00:01:05.66" heatid="36003" lane="3" />
                <ENTRY eventid="38" entrytime="00:02:07.74" heatid="38002" lane="2" />
                <ENTRY eventid="16" entrytime="00:00:59.30" heatid="16001" lane="3" />
                <ENTRY eventid="50" entrytime="00:01:09.55" heatid="50001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="364" eventid="2" swimtime="00:00:59.30" lane="5" heatid="2004" points="579" />
                <RESULT resultid="365" eventid="8" swimtime="00:02:22.61" lane="3" heatid="8002" points="483">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="828" eventid="16" swimtime="00:00:59.18" lane="3" heatid="16001" points="583" />
                <RESULT resultid="366" eventid="24" swimtime="00:02:23.58" lane="8" heatid="24004" points="500">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="367" eventid="28" swimtime="00:00:27.13" lane="7" heatid="28006" points="553" />
                <RESULT resultid="368" eventid="36" swimtime="00:01:09.55" lane="3" heatid="36003" points="408" />
                <RESULT resultid="369" eventid="38" swimtime="00:02:14.77" lane="2" heatid="38002" points="548">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="916" eventid="50" swimtime="00:01:05.80" lane="8" heatid="50001" points="482" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="77" birthdate="2014-01-01" gender="M" lastname="Salfitzky" firstname="Benno" license="448061" nation="GER">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:02:37.53" heatid="8002" lane="2" />
                <ENTRY eventid="12" entrytime="00:01:08.67" heatid="12002" lane="8" />
                <ENTRY eventid="22" entrytime="00:00:34.90" heatid="22002" lane="5" />
                <ENTRY eventid="28" entrytime="00:00:32.87" heatid="28003" lane="2" />
                <ENTRY eventid="36" entrytime="00:01:14.92" heatid="36003" lane="1" />
                <ENTRY eventid="40" entrytime="00:00:30.01" heatid="40002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="370" eventid="8" swimtime="00:02:42.26" lane="2" heatid="8002" points="328">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="371" eventid="12" swimtime="00:01:07.55" lane="8" heatid="12002" points="324" />
                <RESULT resultid="372" eventid="22" swimtime="00:00:34.60" lane="5" heatid="22002" points="315" />
                <RESULT resultid="373" eventid="28" swimtime="00:00:33.12" lane="2" heatid="28003" points="304" />
                <RESULT resultid="374" eventid="36" swimtime="00:01:16.10" lane="1" heatid="36003" points="311" />
                <RESULT resultid="375" eventid="40" swimtime="00:00:29.71" lane="4" heatid="40002" points="348" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="78" birthdate="2012-01-01" gender="M" lastname="Kolkowski" firstname="Daniel" license="443040" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:10:05.22" heatid="10001" lane="5" />
                <ENTRY eventid="22" entrytime="00:00:32.97" heatid="22003" lane="8" />
                <ENTRY eventid="28" entrytime="00:00:30.53" heatid="28004" lane="2" />
                <ENTRY eventid="40" entrytime="00:00:30.18" heatid="40002" lane="5" />
                <ENTRY eventid="46" entrytime="00:04:49.53" heatid="46000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="376" eventid="10" swimtime="00:10:02.72" lane="5" heatid="10001" points="422">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="200" swimtime="00:02:21.81" />
                    <SPLIT distance="300" swimtime="00:03:38.11" />
                    <SPLIT distance="400" swimtime="00:04:54.59" />
                    <SPLIT distance="500" swimtime="00:06:11.45" />
                    <SPLIT distance="600" swimtime="00:07:29.08" />
                    <SPLIT distance="700" swimtime="00:08:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="377" eventid="22" swimtime="00:00:33.33" lane="8" heatid="22003" points="352" />
                <RESULT resultid="378" eventid="28" swimtime="00:00:31.49" lane="2" heatid="28004" points="353" />
                <RESULT resultid="379" eventid="40" status="WDR" swimtime="00:00:00.00" lane="5" heatid="40002" />
                <RESULT resultid="380" eventid="46" status="WDR" swimtime="00:00:00.00" lane="0" heatid="46000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="79" birthdate="2014-01-01" gender="M" lastname="Müller" firstname="Felix" license="447956" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:30.53" heatid="4002" lane="6" />
                <ENTRY eventid="12" entrytime="00:01:08.57" heatid="12002" lane="1" />
                <ENTRY eventid="24" entrytime="00:02:51.88" heatid="24001" lane="4" />
                <ENTRY eventid="30" entrytime="00:03:37.63" heatid="30001" lane="2" />
                <ENTRY eventid="40" entrytime="00:00:30.47" heatid="40002" lane="3" />
                <ENTRY eventid="42" entrytime="00:06:38.84" heatid="42002" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="381" eventid="4" swimtime="00:02:35.17" lane="6" heatid="4002" points="284">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="382" eventid="12" swimtime="00:01:09.32" lane="1" heatid="12002" points="299" />
                <RESULT resultid="383" eventid="24" swimtime="00:02:50.02" lane="4" heatid="24001" points="301">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="384" eventid="30" swimtime="00:03:22.07" lane="2" heatid="30001" points="239">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="385" eventid="40" swimtime="00:00:31.16" lane="3" heatid="40002" points="302" />
                <RESULT resultid="386" eventid="42" swimtime="00:06:00.45" lane="6" heatid="42002" points="304">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.24" />
                    <SPLIT distance="200" swimtime="00:02:56.86" />
                    <SPLIT distance="300" swimtime="00:04:42.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="80" birthdate="2011-01-01" gender="F" lastname="Bürger" firstname="Hannah Victoria" license="424897" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:16.82" heatid="5003" lane="3" />
                <ENTRY eventid="11" entrytime="00:01:01.37" heatid="11003" lane="6" />
                <ENTRY eventid="27" entrytime="00:00:28.62" heatid="27005" lane="5" />
                <ENTRY eventid="35" entrytime="00:01:06.21" heatid="35004" lane="4" />
                <ENTRY eventid="39" entrytime="00:00:28.25" heatid="39004" lane="2" />
                <ENTRY eventid="17" entrytime="00:01:18.73" heatid="17001" lane="3" />
                <ENTRY eventid="31" entrytime="00:01:00.74" heatid="31001" lane="4" />
                <ENTRY eventid="47" entrytime="00:01:08.38" heatid="47001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="387" eventid="5" swimtime="00:01:18.73" lane="3" heatid="5003" points="540" />
                <RESULT resultid="388" eventid="11" swimtime="00:01:00.74" lane="6" heatid="11003" points="617" />
                <RESULT resultid="835" eventid="17" swimtime="00:01:17.79" lane="3" heatid="17001" points="560" />
                <RESULT resultid="389" eventid="27" swimtime="00:00:29.24" lane="5" heatid="27005" points="583" />
                <RESULT resultid="856" eventid="31" swimtime="00:01:00.94" lane="4" heatid="31001" points="610" />
                <RESULT resultid="390" eventid="35" swimtime="00:01:08.38" lane="4" heatid="35004" points="583" />
                <RESULT resultid="391" eventid="39" swimtime="00:00:28.65" lane="2" heatid="39004" points="559" />
                <RESULT resultid="888" eventid="47" swimtime="00:01:07.10" lane="4" heatid="47001" points="617" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="81" birthdate="2008-01-01" gender="F" lastname="Göde" firstname="Helena" license="391855" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:03.80" heatid="1002" lane="4" />
                <ENTRY eventid="11" entrytime="00:00:58.63" heatid="11004" lane="4" />
                <ENTRY eventid="35" entrytime="00:01:09.91" heatid="35005" lane="6" />
                <ENTRY eventid="39" entrytime="00:00:27.27" heatid="39005" lane="2" />
                <ENTRY eventid="14" entrytime="00:01:06.06" heatid="14001" lane="5" />
                <ENTRY eventid="32" entrytime="00:01:00.54" heatid="32001" lane="6" />
                <ENTRY eventid="48" entrytime="00:01:09.73" heatid="48001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="392" eventid="1" swimtime="00:01:06.06" lane="4" heatid="1002" points="582" />
                <RESULT resultid="393" eventid="11" swimtime="00:01:00.54" lane="4" heatid="11004" points="623" />
                <RESULT resultid="814" eventid="14" swimtime="00:01:05.84" lane="5" heatid="14001" points="588" />
                <RESULT resultid="867" eventid="32" swimtime="00:01:00.16" lane="6" heatid="32001" points="635" />
                <RESULT resultid="394" eventid="35" swimtime="00:01:09.73" lane="6" heatid="35005" points="549" />
                <RESULT resultid="395" eventid="39" swimtime="00:00:28.56" lane="2" heatid="39005" points="564" />
                <RESULT resultid="898" eventid="48" swimtime="00:01:09.41" lane="3" heatid="48001" points="557" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="82" birthdate="2012-01-01" gender="F" lastname="Kobus" firstname="Henrijette" license="439567" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:11.61" heatid="1004" lane="7" />
                <ENTRY eventid="23" entrytime="00:02:33.83" heatid="23004" lane="6" />
                <ENTRY eventid="27" entrytime="00:00:31.22" heatid="27004" lane="8" />
                <ENTRY eventid="35" entrytime="00:01:10.18" heatid="35003" lane="6" />
                <ENTRY eventid="39" entrytime="00:00:28.26" heatid="39004" lane="7" />
                <ENTRY eventid="47" entrytime="00:01:11.78" heatid="47001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="396" eventid="1" swimtime="00:01:11.87" lane="7" heatid="1004" points="452" />
                <RESULT resultid="397" eventid="23" swimtime="00:02:38.12" lane="6" heatid="23004" points="507">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="398" eventid="27" swimtime="00:00:30.96" lane="8" heatid="27004" points="491" />
                <RESULT resultid="399" eventid="35" swimtime="00:01:11.78" lane="6" heatid="35003" points="504" />
                <RESULT resultid="400" eventid="39" swimtime="00:00:28.65" lane="7" heatid="39004" points="559" />
                <RESULT resultid="894" eventid="47" swimtime="00:01:11.55" lane="1" heatid="47001" points="509" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="83" birthdate="2008-01-01" gender="M" lastname="Silex" firstname="Konstantin" license="387209" nation="GER">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:02:05.83" heatid="8003" lane="3" />
                <ENTRY eventid="24" entrytime="00:02:14.80" heatid="24004" lane="6" />
                <ENTRY eventid="36" entrytime="00:00:59.27" heatid="36004" lane="5" />
                <ENTRY eventid="44" entrytime="00:00:31.08" heatid="44003" lane="6" />
                <ENTRY eventid="50" entrytime="00:01:01.47" heatid="50001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="401" eventid="8" swimtime="00:02:12.21" lane="3" heatid="8003" points="606">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="402" eventid="24" swimtime="00:02:15.47" lane="6" heatid="24004" points="595">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="403" eventid="36" swimtime="00:01:01.47" lane="5" heatid="36004" points="591" />
                <RESULT resultid="404" eventid="44" swimtime="00:00:32.52" lane="6" heatid="44003" points="508" />
                <RESULT resultid="910" eventid="50" swimtime="00:01:01.31" lane="5" heatid="50001" points="596" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="84" birthdate="2011-01-01" gender="F" lastname="Winkler" firstname="Maike" license="424911" nation="GER">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:01:00.69" heatid="11004" lane="3" />
                <ENTRY eventid="23" entrytime="00:02:28.81" heatid="23005" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:29.21" heatid="27005" lane="6" />
                <ENTRY eventid="39" entrytime="00:00:27.05" heatid="39005" lane="3" />
                <ENTRY eventid="45" entrytime="00:04:46.48" heatid="45003" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:01.36" heatid="31001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="405" eventid="11" swimtime="00:01:01.36" lane="3" heatid="11004" points="598" />
                <RESULT resultid="406" eventid="23" swimtime="00:02:34.39" lane="1" heatid="23005" points="545">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="407" eventid="27" swimtime="00:00:29.25" lane="6" heatid="27005" points="582" />
                <RESULT resultid="859" eventid="31" swimtime="00:01:02.18" lane="6" heatid="31001" points="575" />
                <RESULT resultid="408" eventid="39" swimtime="00:00:27.78" lane="3" heatid="39005" points="613" />
                <RESULT resultid="409" eventid="45" swimtime="00:04:48.46" lane="4" heatid="45003" points="543">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.81" />
                    <SPLIT distance="200" swimtime="00:02:20.04" />
                    <SPLIT distance="300" swimtime="00:03:34.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="85" birthdate="2012-01-01" gender="M" lastname="Martin" firstname="Mika-Frederik" license="436899" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:03.01" heatid="2003" lane="3" />
                <ENTRY eventid="6" entrytime="00:01:17.42" heatid="6003" lane="3" />
                <ENTRY eventid="22" entrytime="00:00:31.82" heatid="22003" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:27.14" heatid="28006" lane="1" />
                <ENTRY eventid="15" entrytime="00:01:02.15" heatid="15001" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:15.93" heatid="19001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="410" eventid="2" swimtime="00:01:02.15" lane="3" heatid="2003" points="503" />
                <RESULT resultid="411" eventid="6" swimtime="00:01:15.93" lane="3" heatid="6003" points="420" />
                <RESULT resultid="818" eventid="15" swimtime="00:01:03.23" lane="4" heatid="15001" points="478" />
                <RESULT resultid="849" eventid="19" swimtime="00:01:19.59" lane="2" heatid="19001" points="365" />
                <RESULT resultid="412" eventid="22" swimtime="00:00:33.13" lane="1" heatid="22003" points="359" />
                <RESULT resultid="413" eventid="28" swimtime="00:00:28.18" lane="1" heatid="28006" points="493" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="86" birthdate="2011-01-01" gender="F" lastname="Mauermann" firstname="Mila" license="424568" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:05.65" heatid="1003" lane="3" />
                <ENTRY eventid="11" entrytime="00:01:00.89" heatid="11003" lane="3" />
                <ENTRY eventid="23" entrytime="00:02:28.78" heatid="23005" lane="7" />
                <ENTRY eventid="35" entrytime="00:01:10.77" heatid="35005" lane="2" />
                <ENTRY eventid="39" entrytime="00:00:28.02" heatid="39004" lane="6" />
                <ENTRY eventid="13" entrytime="00:01:09.13" heatid="13001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="414" eventid="1" swimtime="00:01:09.13" lane="3" heatid="1003" points="508" />
                <RESULT resultid="415" eventid="11" swimtime="00:01:03.76" lane="3" heatid="11003" points="533" />
                <RESULT resultid="804" eventid="13" swimtime="00:01:08.51" lane="5" heatid="13001" points="522" />
                <RESULT resultid="416" eventid="23" swimtime="00:02:35.70" lane="7" heatid="23005" points="531">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="417" eventid="35" swimtime="00:01:13.65" lane="2" heatid="35005" points="466" />
                <RESULT resultid="418" eventid="39" swimtime="00:00:29.15" lane="6" heatid="39004" points="531" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="87" birthdate="2013-01-01" gender="M" lastname="Wiese" firstname="Niklas" license="445789" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:10:43.87" heatid="10001" lane="2" />
                <ENTRY eventid="24" entrytime="00:02:44.95" heatid="24002" lane="8" />
                <ENTRY eventid="28" entrytime="00:00:36.25" heatid="28002" lane="2" />
                <ENTRY eventid="40" entrytime="00:00:33.54" heatid="40001" lane="2" />
                <ENTRY eventid="46" entrytime="00:05:07.14" heatid="46002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="419" eventid="10" swimtime="00:10:38.82" lane="2" heatid="10001" points="354">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="200" swimtime="00:02:32.65" />
                    <SPLIT distance="300" swimtime="00:03:53.27" />
                    <SPLIT distance="400" swimtime="00:05:14.76" />
                    <SPLIT distance="500" swimtime="00:06:37.27" />
                    <SPLIT distance="600" swimtime="00:07:59.46" />
                    <SPLIT distance="700" swimtime="00:09:20.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="420" eventid="24" swimtime="00:02:43.91" lane="8" heatid="24002" points="336">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="421" eventid="28" swimtime="00:00:36.36" lane="2" heatid="28002" points="229" />
                <RESULT resultid="422" eventid="40" swimtime="00:00:33.35" lane="2" heatid="40001" points="246" />
                <RESULT resultid="423" eventid="46" swimtime="00:05:13.37" lane="1" heatid="46002" points="346">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="200" swimtime="00:02:34.71" />
                    <SPLIT distance="300" swimtime="00:03:55.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="88" birthdate="2013-01-01" gender="M" lastname="Gruhl" firstname="Theodor" license="445434" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:28.65" heatid="6001" lane="6" />
                <ENTRY eventid="8" entrytime="00:02:55.64" heatid="8001" lane="5" />
                <ENTRY eventid="22" entrytime="00:00:37.88" heatid="22002" lane="1" />
                <ENTRY eventid="30" entrytime="00:03:09.87" heatid="30001" lane="6" />
                <ENTRY eventid="36" entrytime="00:01:21.08" heatid="36001" lane="3" />
                <ENTRY eventid="40" entrytime="00:00:32.38" heatid="40001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="424" eventid="6" swimtime="00:01:30.14" lane="6" heatid="6001" points="251" />
                <RESULT resultid="425" eventid="8" swimtime="00:02:58.48" lane="5" heatid="8001" points="246">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="426" eventid="22" swimtime="00:00:37.92" lane="1" heatid="22002" points="239" />
                <RESULT resultid="427" eventid="30" swimtime="00:03:07.34" lane="6" heatid="30001" points="300">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="428" eventid="36" swimtime="00:01:24.33" lane="3" heatid="36001" points="229" />
                <RESULT resultid="429" eventid="40" swimtime="00:00:31.66" lane="5" heatid="40001" points="288" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Landesschwimmverband Sachsen-Anhalt" nation="GER" region="13" code="13">
          <ATHLETES>
            <ATHLETE athleteid="170" birthdate="2012-01-01" gender="M" lastname="Tietje" firstname="Fabian" license="434342" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:00:00.00" heatid="4002" lane="8" />
                <ENTRY eventid="24" entrytime="00:00:00.00" heatid="24004" lane="4" />
                <ENTRY eventid="8" entrytime="00:00:00.00" heatid="8002" lane="1" />
                <ENTRY eventid="36" entrytime="00:00:00.00" heatid="36001" lane="1" />
                <ENTRY eventid="46" entrytime="00:00:00.00" heatid="46001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="798" eventid="4" swimtime="00:02:24.15" lane="8" heatid="4002" points="354">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="800" eventid="8" swimtime="00:02:39.51" lane="1" heatid="8002" points="345">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="799" eventid="24" status="DSQ" swimtime="00:02:40.37" lane="4" heatid="24004" comment="Sportler startete vor dem Startsignal.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="801" eventid="36" swimtime="00:01:10.77" lane="1" heatid="36001" points="387" />
                <RESULT resultid="802" eventid="46" swimtime="00:05:07.50" lane="2" heatid="46001" points="366">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="200" swimtime="00:02:28.90" />
                    <SPLIT distance="300" swimtime="00:03:49.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Chemnitz von 1892" nation="GER" region="12" code="3353">
          <ATHLETES>
            <ATHLETE athleteid="49" birthdate="2005-01-01" gender="M" lastname="Rèvèsz" firstname="Enzio" license="325104" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:01:54.85" heatid="4004" lane="5" />
                <ENTRY eventid="24" entrytime="00:02:06.38" heatid="24004" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="242" eventid="4" swimtime="00:01:55.07" lane="5" heatid="4004" points="696">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="243" eventid="24" swimtime="00:02:10.74" lane="5" heatid="24004" points="662">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="50" birthdate="2009-01-01" gender="M" lastname="Seidel" firstname="Gustav" license="365674" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:08.39" heatid="4003" lane="2" />
                <ENTRY eventid="10" entrytime="00:09:06.86" heatid="10002" lane="3" />
                <ENTRY eventid="22" entrytime="00:00:30.66" heatid="22003" lane="7" />
                <ENTRY eventid="36" entrytime="00:01:05.99" heatid="36004" lane="6" />
                <ENTRY eventid="46" entrytime="00:04:25.39" heatid="46003" lane="2" />
                <ENTRY eventid="50" entrytime="00:01:06.32" heatid="50001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="244" eventid="4" swimtime="00:02:10.17" lane="2" heatid="4003" points="481">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="245" eventid="10" swimtime="00:09:23.97" lane="3" heatid="10002" points="515">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.31" />
                    <SPLIT distance="200" swimtime="00:02:16.59" />
                    <SPLIT distance="300" swimtime="00:03:27.28" />
                    <SPLIT distance="400" swimtime="00:04:38.48" />
                    <SPLIT distance="500" swimtime="00:05:49.92" />
                    <SPLIT distance="600" swimtime="00:07:01.90" />
                    <SPLIT distance="700" swimtime="00:08:14.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="246" eventid="22" swimtime="00:00:30.73" lane="7" heatid="22003" points="450" />
                <RESULT resultid="247" eventid="36" swimtime="00:01:06.32" lane="6" heatid="36004" points="470" />
                <RESULT resultid="248" eventid="46" swimtime="00:04:35.17" lane="2" heatid="46003" points="511">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="200" swimtime="00:02:14.65" />
                    <SPLIT distance="300" swimtime="00:03:25.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="913" eventid="50" swimtime="00:01:06.62" lane="2" heatid="50001" points="464" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="51" birthdate="2011-01-01" gender="F" lastname="Schultze" firstname="Heidi" license="423424" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:14.18" heatid="1004" lane="8" />
                <ENTRY eventid="7" entrytime="00:02:44.17" heatid="7001" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:42.85" heatid="23003" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:33.87" heatid="27003" lane="8" />
                <ENTRY eventid="35" entrytime="00:01:19.75" heatid="35002" lane="2" />
                <ENTRY eventid="45" entrytime="00:05:03.76" heatid="45003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="249" eventid="1" swimtime="00:01:16.85" lane="8" heatid="1004" points="370" />
                <RESULT resultid="250" eventid="7" swimtime="00:02:42.30" lane="5" heatid="7001" points="436">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="251" eventid="23" swimtime="00:02:43.86" lane="2" heatid="23003" points="455">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="252" eventid="27" swimtime="00:00:34.11" lane="8" heatid="27003" points="367" />
                <RESULT resultid="253" eventid="35" swimtime="00:01:17.24" lane="2" heatid="35002" points="404" />
                <RESULT resultid="254" eventid="45" swimtime="00:05:14.49" lane="2" heatid="45003" points="419">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                    <SPLIT distance="200" swimtime="00:02:32.61" />
                    <SPLIT distance="300" swimtime="00:03:54.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="52" birthdate="2010-01-01" gender="M" lastname="Postel" firstname="Jannek" license="408981" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:13.01" heatid="6002" lane="5" />
                <ENTRY eventid="12" entrytime="00:00:59.96" heatid="12004" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:30.63" heatid="28004" lane="7" />
                <ENTRY eventid="36" entrytime="00:01:08.77" heatid="36003" lane="2" />
                <ENTRY eventid="44" entrytime="00:00:32.32" heatid="44003" lane="2" />
                <ENTRY eventid="19" entrytime="00:01:10.66" heatid="19001" lane="4" />
                <ENTRY eventid="33" entrytime="00:00:59.12" heatid="33001" lane="2" />
                <ENTRY eventid="49" entrytime="00:01:06.49" heatid="49001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="255" eventid="6" swimtime="00:01:10.66" lane="5" heatid="6002" points="521" />
                <RESULT resultid="256" eventid="12" swimtime="00:00:59.12" lane="1" heatid="12004" points="483" />
                <RESULT resultid="845" eventid="19" swimtime="00:01:09.64" lane="4" heatid="19001" points="544" />
                <RESULT resultid="257" eventid="28" swimtime="00:00:28.29" lane="7" heatid="28004" points="487" />
                <RESULT resultid="875" eventid="33" swimtime="00:00:59.03" lane="2" heatid="33001" points="485" />
                <RESULT resultid="258" eventid="36" swimtime="00:01:06.49" lane="2" heatid="36003" points="467" />
                <RESULT resultid="259" eventid="44" swimtime="00:00:32.96" lane="2" heatid="44003" points="488" />
                <RESULT resultid="902" eventid="49" swimtime="00:01:05.94" lane="5" heatid="49001" points="479" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="53" birthdate="2008-01-01" gender="F" lastname="Bergmann" firstname="Kristin" license="364361" nation="GER">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:00:59.45" heatid="11005" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:23.90" heatid="23005" lane="3" />
                <ENTRY eventid="35" entrytime="00:01:05.81" heatid="35005" lane="4" />
                <ENTRY eventid="39" entrytime="00:00:27.28" heatid="39005" lane="7" />
                <ENTRY eventid="32" entrytime="00:00:58.95" heatid="32001" lane="5" />
                <ENTRY eventid="48" entrytime="00:01:06.97" heatid="48001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="260" eventid="11" swimtime="00:00:58.95" lane="5" heatid="11005" points="674" />
                <RESULT resultid="261" eventid="23" swimtime="00:02:23.74" lane="3" heatid="23005" points="675">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="865" eventid="32" swimtime="00:00:58.82" lane="5" heatid="32001" points="679" />
                <RESULT resultid="262" eventid="35" swimtime="00:01:06.97" lane="4" heatid="35005" points="620" />
                <RESULT resultid="263" eventid="39" swimtime="00:00:27.75" lane="7" heatid="39005" points="615" />
                <RESULT resultid="896" eventid="48" swimtime="00:01:07.32" lane="4" heatid="48001" points="611" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="54" birthdate="2010-01-01" gender="F" lastname="Ahnert" firstname="Lina Jolie" license="410263" nation="GER">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:02:32.66" heatid="7002" lane="3" />
                <ENTRY eventid="21" entrytime="00:00:32.04" heatid="21003" lane="6" />
                <ENTRY eventid="35" entrytime="00:01:08.49" heatid="35004" lane="5" />
                <ENTRY eventid="39" entrytime="00:00:29.38" heatid="39003" lane="7" />
                <ENTRY eventid="47" entrytime="00:01:10.58" heatid="47001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="264" eventid="7" swimtime="00:02:33.72" lane="3" heatid="7002" points="514">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="265" eventid="21" swimtime="00:00:32.58" lane="6" heatid="21003" points="560" />
                <RESULT resultid="266" eventid="35" swimtime="00:01:10.58" lane="5" heatid="35004" points="530" />
                <RESULT resultid="267" eventid="39" status="DNS" swimtime="00:00:00.00" lane="7" heatid="39003" />
                <RESULT resultid="891" eventid="47" swimtime="00:01:11.75" lane="6" heatid="47001" points="504" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="55" birthdate="2011-01-01" gender="F" lastname="Franke" firstname="Loreley" license="447682" nation="GER">
              <ENTRIES>
                <ENTRY eventid="11" entrytime="00:01:05.92" heatid="11005" lane="8" />
                <ENTRY eventid="23" entrytime="00:02:44.18" heatid="23002" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:31.86" heatid="27003" lane="5" />
                <ENTRY eventid="35" entrytime="00:01:16.82" heatid="35002" lane="5" />
                <ENTRY eventid="39" entrytime="00:00:29.57" heatid="39003" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="268" eventid="11" swimtime="00:01:05.77" lane="8" heatid="11005" points="486" />
                <RESULT resultid="269" eventid="23" swimtime="00:02:41.60" lane="4" heatid="23002" points="475">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="270" eventid="27" swimtime="00:00:31.34" lane="5" heatid="27003" points="473" />
                <RESULT resultid="271" eventid="35" swimtime="00:01:15.13" lane="5" heatid="35002" points="439" />
                <RESULT resultid="272" eventid="39" swimtime="00:00:29.98" lane="8" heatid="39003" points="488" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="56" birthdate="2007-01-01" gender="M" lastname="Seifert" firstname="Luca" license="370516" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:01.12" heatid="4004" lane="1" />
                <ENTRY eventid="12" entrytime="00:00:56.28" heatid="12004" lane="6" />
                <ENTRY eventid="22" entrytime="00:00:26.90" heatid="22003" lane="4" />
                <ENTRY eventid="36" entrytime="00:00:57.84" heatid="36003" lane="4" />
                <ENTRY eventid="40" entrytime="00:00:25.72" heatid="40005" lane="1" />
                <ENTRY eventid="34" entrytime="00:00:55.19" heatid="34001" lane="1" />
                <ENTRY eventid="50" entrytime="00:00:58.57" heatid="50001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="273" eventid="4" swimtime="00:02:00.87" lane="1" heatid="4004" points="600">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="274" eventid="12" swimtime="00:00:55.19" lane="6" heatid="12004" points="594" />
                <RESULT resultid="275" eventid="22" swimtime="00:00:27.35" lane="4" heatid="22003" points="638" />
                <RESULT resultid="886" eventid="34" swimtime="00:00:54.98" lane="1" heatid="34001" points="601" />
                <RESULT resultid="276" eventid="36" swimtime="00:00:58.57" lane="4" heatid="36003" points="683" />
                <RESULT resultid="277" eventid="40" swimtime="00:00:25.70" lane="1" heatid="40005" points="538" />
                <RESULT resultid="909" eventid="50" swimtime="00:00:58.50" lane="4" heatid="50001" points="686" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="57" birthdate="2006-01-01" gender="M" lastname="Bergmann" firstname="Magnus" license="352440" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:01:53.44" heatid="4004" lane="4" />
                <ENTRY eventid="12" entrytime="00:00:53.21" heatid="12005" lane="4" />
                <ENTRY eventid="46" entrytime="00:03:59.96" heatid="46003" lane="4" />
                <ENTRY eventid="34" entrytime="00:00:54.11" heatid="34001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="278" eventid="4" swimtime="00:01:55.00" lane="4" heatid="4004" points="697">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="279" eventid="12" swimtime="00:00:54.11" lane="4" heatid="12005" points="630" />
                <RESULT resultid="881" eventid="34" swimtime="00:00:53.80" lane="5" heatid="34001" points="641" />
                <RESULT resultid="280" eventid="46" swimtime="00:04:04.67" lane="4" heatid="46003" points="727">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.28" />
                    <SPLIT distance="200" swimtime="00:01:59.09" />
                    <SPLIT distance="300" swimtime="00:03:02.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="58" birthdate="2011-01-01" gender="F" lastname="Schreiber" firstname="Marlene" license="423429">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:18.39" heatid="3002" lane="3" />
                <ENTRY eventid="21" entrytime="00:00:30.48" heatid="21003" lane="4" />
                <ENTRY eventid="37" entrytime="00:02:56.31" heatid="37002" lane="1" />
                <ENTRY eventid="43" entrytime="00:00:38.34" heatid="43002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="281" eventid="3" swimtime="00:02:15.00" lane="3" heatid="3002" points="574">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="282" eventid="21" swimtime="00:00:31.98" lane="4" heatid="21003" points="592" />
                <RESULT resultid="283" eventid="37" swimtime="00:02:41.85" lane="1" heatid="37002" points="426">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="284" eventid="43" swimtime="00:00:36.46" lane="4" heatid="43002" points="511" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="59" birthdate="2009-01-01" gender="F" lastname="Nitschke" firstname="Melina" license="391097" nation="GER">
              <ENTRIES>
                <ENTRY eventid="9" entrytime="00:09:03.21" heatid="9002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="285" eventid="9" swimtime="00:09:03.74" lane="4" heatid="9002" points="708">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.53" />
                    <SPLIT distance="200" swimtime="00:02:10.60" />
                    <SPLIT distance="300" swimtime="00:03:18.40" />
                    <SPLIT distance="400" swimtime="00:04:26.53" />
                    <SPLIT distance="500" swimtime="00:05:35.13" />
                    <SPLIT distance="600" swimtime="00:06:44.39" />
                    <SPLIT distance="700" swimtime="00:07:54.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="60" birthdate="2010-01-01" gender="F" lastname="Naumann" firstname="Noelle" license="408977" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:14.21" heatid="3002" lane="4" />
                <ENTRY eventid="7" entrytime="00:02:34.55" heatid="7002" lane="1" />
                <ENTRY eventid="21" entrytime="00:00:34.39" heatid="21002" lane="5" />
                <ENTRY eventid="35" entrytime="00:01:13.57" heatid="35005" lane="1" />
                <ENTRY eventid="39" entrytime="00:00:28.38" heatid="39004" lane="1" />
                <ENTRY eventid="47" entrytime="00:01:11.79" heatid="47001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="286" eventid="3" swimtime="00:02:14.23" lane="4" heatid="3002" points="584">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="287" eventid="7" swimtime="00:02:34.91" lane="1" heatid="7002" points="502">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="288" eventid="21" swimtime="00:00:33.72" lane="5" heatid="21002" points="505" />
                <RESULT resultid="289" eventid="35" swimtime="00:01:11.79" lane="1" heatid="35005" points="503" />
                <RESULT resultid="290" eventid="39" swimtime="00:00:28.21" lane="1" heatid="39004" points="586" />
                <RESULT resultid="895" eventid="47" swimtime="00:01:11.90" lane="8" heatid="47001" points="501" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="61" birthdate="2011-01-01" gender="M" lastname="Wehner" firstname="Paul" license="423422">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:10.74" heatid="2003" lane="1" />
                <ENTRY eventid="12" entrytime="00:01:00.57" heatid="12003" lane="8" />
                <ENTRY eventid="28" entrytime="00:00:31.10" heatid="28004" lane="1" />
                <ENTRY eventid="38" entrytime="00:02:26.71" heatid="38002" lane="1" />
                <ENTRY eventid="42" entrytime="00:05:21.93" heatid="42003" lane="6" />
                <ENTRY eventid="15" entrytime="00:01:05.38" heatid="15001" lane="1" />
                <ENTRY eventid="33" entrytime="00:00:59.80" heatid="33001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="291" eventid="2" swimtime="00:01:05.38" lane="1" heatid="2003" points="432" />
                <RESULT resultid="292" eventid="12" swimtime="00:00:59.80" lane="8" heatid="12003" points="467" />
                <RESULT resultid="824" eventid="15" swimtime="00:01:04.60" lane="1" heatid="15001" points="448" />
                <RESULT resultid="293" eventid="28" swimtime="00:00:30.03" lane="1" heatid="28004" points="407" />
                <RESULT resultid="878" eventid="33" swimtime="00:01:00.13" lane="8" heatid="33001" points="459" />
                <RESULT resultid="294" eventid="38" swimtime="00:02:27.45" lane="1" heatid="38002" points="419">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="295" eventid="42" status="DSQ" swimtime="00:05:26.60" lane="6" heatid="42003" comment="Die Rückenstrecke wurde nicht in Rückenlage beendet.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="200" swimtime="00:02:41.18" />
                    <SPLIT distance="300" swimtime="00:04:14.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="62" birthdate="2011-01-01" gender="M" lastname="Stang" firstname="Philipp" license="423425">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:17.21" heatid="4002" lane="5" />
                <ENTRY eventid="12" entrytime="00:01:05.01" heatid="12002" lane="6" />
                <ENTRY eventid="28" entrytime="00:00:32.57" heatid="28003" lane="3" />
                <ENTRY eventid="40" entrytime="00:00:29.89" heatid="40003" lane="1" />
                <ENTRY eventid="46" entrytime="00:04:42.89" heatid="46003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="296" eventid="4" swimtime="00:02:17.25" lane="5" heatid="4002" points="410">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="297" eventid="12" swimtime="00:01:04.08" lane="6" heatid="12002" points="379" />
                <RESULT resultid="298" eventid="28" swimtime="00:00:31.88" lane="3" heatid="28003" points="340" />
                <RESULT resultid="299" eventid="40" swimtime="00:00:29.38" lane="1" heatid="40003" points="360" />
                <RESULT resultid="300" eventid="46" swimtime="00:04:44.79" lane="1" heatid="46003" points="461">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                    <SPLIT distance="200" swimtime="00:02:20.29" />
                    <SPLIT distance="300" swimtime="00:03:33.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="63" birthdate="2012-01-01" gender="F" lastname="Drechsel" firstname="Rosalie" license="437426" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:12.70" heatid="1002" lane="7" />
                <ENTRY eventid="11" entrytime="00:01:07.38" heatid="11003" lane="8" />
                <ENTRY eventid="23" entrytime="00:02:40.27" heatid="23003" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:33.27" heatid="27003" lane="7" />
                <ENTRY eventid="41" entrytime="00:05:37.91" heatid="41000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="301" eventid="1" status="WDR" swimtime="00:00:00.00" lane="7" heatid="1002" />
                <RESULT resultid="302" eventid="11" status="WDR" swimtime="00:00:00.00" lane="8" heatid="11003" />
                <RESULT resultid="303" eventid="23" status="WDR" swimtime="00:00:00.00" lane="3" heatid="23003" />
                <RESULT resultid="304" eventid="27" status="WDR" swimtime="00:00:00.00" lane="7" heatid="27003" />
                <RESULT resultid="305" eventid="41" status="WDR" swimtime="00:00:00.00" lane="0" heatid="41000" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC DHfK Leipzig" nation="GER" region="12" code="3354">
          <ATHLETES>
            <ATHLETE athleteid="4" birthdate="2011-01-01" gender="M" lastname="Milbach" firstname="Mio Moritz" license="408265" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:22.36" heatid="2002" lane="2" />
                <ENTRY eventid="6" entrytime="00:01:32.25" heatid="6001" lane="2" />
                <ENTRY eventid="24" entrytime="00:02:44.59" heatid="24002" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:35.37" heatid="28002" lane="3" />
                <ENTRY eventid="36" entrytime="00:01:16.31" heatid="36002" lane="1" />
                <ENTRY eventid="44" entrytime="00:00:40.64" heatid="44002" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="12" eventid="2" swimtime="00:01:20.90" lane="2" heatid="2002" points="228" />
                <RESULT resultid="13" eventid="6" swimtime="00:01:27.06" lane="2" heatid="6001" points="278" />
                <RESULT resultid="14" eventid="24" swimtime="00:02:46.33" lane="1" heatid="24002" points="321">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="15" eventid="28" swimtime="00:00:35.26" lane="3" heatid="28002" points="251" />
                <RESULT resultid="16" eventid="36" swimtime="00:01:18.16" lane="1" heatid="36002" points="287" />
                <RESULT resultid="17" eventid="44" swimtime="00:00:40.41" lane="7" heatid="44002" points="264" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Freital" nation="GER" region="12" code="3339">
          <ATHLETES>
            <ATHLETE athleteid="5" birthdate="2009-01-01" gender="F" lastname="Lange" firstname="Alia" license="402584">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:02:34.07" heatid="7002" lane="6" />
                <ENTRY eventid="21" entrytime="00:00:32.81" heatid="21003" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:30.44" heatid="27004" lane="5" />
                <ENTRY eventid="39" entrytime="00:00:27.23" heatid="39005" lane="6" />
                <ENTRY eventid="43" entrytime="00:00:39.52" heatid="43002" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="18" eventid="7" swimtime="00:02:32.84" lane="6" heatid="7002" points="522">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="19" eventid="21" swimtime="00:00:33.50" lane="1" heatid="21003" points="515" />
                <RESULT resultid="20" eventid="27" swimtime="00:00:29.78" lane="5" heatid="27004" points="552" />
                <RESULT resultid="21" eventid="39" swimtime="00:00:27.70" lane="6" heatid="39005" points="619" />
                <RESULT resultid="22" eventid="43" swimtime="00:00:37.55" lane="6" heatid="43002" points="468" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="6" birthdate="2011-01-01" gender="F" lastname="Jang" firstname="Jule" license="425575">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:09.30" heatid="1002" lane="6" />
                <ENTRY eventid="5" entrytime="00:01:16.35" heatid="5002" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:31.77" heatid="23004" lane="5" />
                <ENTRY eventid="27" entrytime="00:00:30.83" heatid="27004" lane="3" />
                <ENTRY eventid="35" entrytime="00:01:13.91" heatid="35004" lane="1" />
                <ENTRY eventid="39" entrytime="00:00:27.50" heatid="39004" lane="4" />
                <ENTRY eventid="13" entrytime="00:01:10.06" heatid="13001" lane="6" />
                <ENTRY eventid="17" entrytime="00:01:19.55" heatid="17001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="23" eventid="1" swimtime="00:01:10.06" lane="6" heatid="1002" points="488" />
                <RESULT resultid="24" eventid="5" swimtime="00:01:19.55" lane="5" heatid="5002" points="523" />
                <RESULT resultid="806" eventid="13" swimtime="00:01:08.39" lane="6" heatid="13001" points="525" />
                <RESULT resultid="837" eventid="17" swimtime="00:01:19.31" lane="2" heatid="17001" points="528" />
                <RESULT resultid="25" eventid="23" swimtime="00:02:32.22" lane="5" heatid="23004" points="568">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="26" eventid="27" swimtime="00:00:30.94" lane="3" heatid="27004" points="492" />
                <RESULT resultid="27" eventid="35" swimtime="00:01:14.71" lane="1" heatid="35004" points="447" />
                <RESULT resultid="28" eventid="39" swimtime="00:00:28.29" lane="4" heatid="39004" points="581" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="7" birthdate="2013-01-01" gender="M" lastname="Tetzlaff" firstname="Luis Max" license="445646">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:10:45.86" heatid="10001" lane="7" />
                <ENTRY eventid="24" entrytime="00:02:41.90" heatid="24002" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:35.35" heatid="28002" lane="5" />
                <ENTRY eventid="40" entrytime="00:00:31.28" heatid="40002" lane="7" />
                <ENTRY eventid="46" entrytime="00:05:05.63" heatid="46002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="29" eventid="10" swimtime="00:10:36.55" lane="7" heatid="10001" points="358">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="200" swimtime="00:02:31.40" />
                    <SPLIT distance="300" swimtime="00:03:53.29" />
                    <SPLIT distance="400" swimtime="00:05:14.93" />
                    <SPLIT distance="500" swimtime="00:06:36.29" />
                    <SPLIT distance="600" swimtime="00:07:57.43" />
                    <SPLIT distance="700" swimtime="00:09:18.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="30" eventid="24" swimtime="00:02:42.07" lane="2" heatid="24002" points="348">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="31" eventid="28" swimtime="00:00:33.67" lane="5" heatid="28002" points="289" />
                <RESULT resultid="32" eventid="40" swimtime="00:00:31.14" lane="7" heatid="40002" points="302" />
                <RESULT resultid="33" eventid="46" swimtime="00:05:12.12" lane="2" heatid="46002" points="350">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.75" />
                    <SPLIT distance="200" swimtime="00:02:33.40" />
                    <SPLIT distance="300" swimtime="00:03:53.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="8" birthdate="2007-01-01" gender="M" lastname="Kovács" firstname="Mika" license="362600">
              <ENTRIES>
                <ENTRY eventid="26" entrytime="00:15:56.45" heatid="26002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="34" eventid="26" swimtime="00:16:45.95" lane="4" heatid="26002" points="648">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.77" />
                    <SPLIT distance="200" swimtime="00:02:06.57" />
                    <SPLIT distance="300" swimtime="00:03:13.34" />
                    <SPLIT distance="400" swimtime="00:04:20.40" />
                    <SPLIT distance="500" swimtime="00:05:27.05" />
                    <SPLIT distance="600" swimtime="00:06:34.07" />
                    <SPLIT distance="700" swimtime="00:07:41.50" />
                    <SPLIT distance="800" swimtime="00:08:48.96" />
                    <SPLIT distance="900" swimtime="00:09:56.71" />
                    <SPLIT distance="1000" swimtime="00:11:04.74" />
                    <SPLIT distance="1100" swimtime="00:12:13.41" />
                    <SPLIT distance="1200" swimtime="00:13:21.73" />
                    <SPLIT distance="1300" swimtime="00:14:30.23" />
                    <SPLIT distance="1400" swimtime="00:15:39.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Magdeburg" nation="GER" region="13" code="3580">
          <ATHLETES>
            <ATHLETE athleteid="120" birthdate="2006-01-01" gender="M" lastname="Schubert" firstname="Arne" license="381621" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:00:56.19" heatid="2003" lane="4" />
                <ENTRY eventid="8" entrytime="00:02:03.19" heatid="8003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="561" eventid="2" status="WDR" swimtime="00:00:00.00" lane="4" heatid="2003" />
                <RESULT resultid="562" eventid="8" status="WDR" swimtime="00:00:00.00" lane="4" heatid="8003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121" birthdate="2011-01-01" gender="M" lastname="Kuzmin" firstname="Artemiy" license="426385" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:14.63" heatid="2004" lane="8" />
                <ENTRY eventid="6" entrytime="00:01:19.08" heatid="6001" lane="3" />
                <ENTRY eventid="26" entrytime="00:20:20.20" heatid="26002" lane="6" />
                <ENTRY eventid="38" entrytime="00:02:46.83" heatid="38001" lane="3" />
                <ENTRY eventid="46" entrytime="00:04:51.94" heatid="46002" lane="6" />
                <ENTRY eventid="19" entrytime="00:01:22.55" heatid="19001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="563" eventid="2" swimtime="00:01:15.05" lane="8" heatid="2004" points="286" />
                <RESULT resultid="564" eventid="6" swimtime="00:01:22.55" lane="3" heatid="6001" points="327" />
                <RESULT resultid="851" eventid="19" swimtime="00:01:20.83" lane="1" heatid="19001" points="348" />
                <RESULT resultid="565" eventid="26" swimtime="00:19:05.92" lane="6" heatid="26002" points="438">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                    <SPLIT distance="200" swimtime="00:02:31.21" />
                    <SPLIT distance="300" swimtime="00:03:47.74" />
                    <SPLIT distance="400" swimtime="00:05:04.67" />
                    <SPLIT distance="500" swimtime="00:06:22.12" />
                    <SPLIT distance="600" swimtime="00:07:39.17" />
                    <SPLIT distance="700" swimtime="00:08:55.91" />
                    <SPLIT distance="800" swimtime="00:10:13.94" />
                    <SPLIT distance="900" swimtime="00:11:30.75" />
                    <SPLIT distance="1000" swimtime="00:12:47.92" />
                    <SPLIT distance="1100" swimtime="00:14:03.73" />
                    <SPLIT distance="1200" swimtime="00:15:20.16" />
                    <SPLIT distance="1300" swimtime="00:16:36.84" />
                    <SPLIT distance="1400" swimtime="00:17:52.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="566" eventid="38" swimtime="00:02:48.62" lane="3" heatid="38001" points="280">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="567" eventid="46" swimtime="00:04:51.57" lane="6" heatid="46002" points="429">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.25" />
                    <SPLIT distance="200" swimtime="00:02:24.18" />
                    <SPLIT distance="300" swimtime="00:03:38.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122" birthdate="2010-01-01" gender="F" lastname="Haubrich" firstname="Caroline" license="406960" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:17.65" heatid="5001" lane="3" />
                <ENTRY eventid="11" entrytime="00:01:03.08" heatid="11004" lane="7" />
                <ENTRY eventid="29" entrytime="00:02:47.34" heatid="29002" lane="5" />
                <ENTRY eventid="35" entrytime="00:01:14.91" heatid="35005" lane="8" />
                <ENTRY eventid="43" entrytime="00:00:35.35" heatid="43003" lane="6" />
                <ENTRY eventid="17" entrytime="00:01:18.20" heatid="17001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="568" eventid="5" swimtime="00:01:18.20" lane="3" heatid="5001" points="551" />
                <RESULT resultid="569" eventid="11" swimtime="00:01:04.23" lane="7" heatid="11004" points="521" />
                <RESULT resultid="834" eventid="17" swimtime="00:01:18.98" lane="5" heatid="17001" points="535" />
                <RESULT resultid="570" eventid="29" swimtime="00:02:51.55" lane="5" heatid="29002" points="515">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="571" eventid="35" swimtime="00:01:14.34" lane="8" heatid="35005" points="453" />
                <RESULT resultid="572" eventid="43" swimtime="00:00:35.89" lane="6" heatid="43003" points="536" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123" birthdate="2014-01-01" gender="M" lastname="Zimmermann" firstname="Claas" license="459680" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:20.48" heatid="2002" lane="3" />
                <ENTRY eventid="12" entrytime="00:01:12.64" heatid="12001" lane="6" />
                <ENTRY eventid="22" entrytime="00:00:36.82" heatid="22002" lane="6" />
                <ENTRY eventid="28" entrytime="00:00:32.56" heatid="28003" lane="5" />
                <ENTRY eventid="40" entrytime="00:00:31.61" heatid="40002" lane="8" />
                <ENTRY eventid="44" entrytime="00:00:46.25" heatid="44001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="573" eventid="2" swimtime="00:01:15.88" lane="3" heatid="2002" points="276" />
                <RESULT resultid="574" eventid="12" swimtime="00:01:12.15" lane="6" heatid="12001" points="265" />
                <RESULT resultid="575" eventid="22" swimtime="00:00:36.27" lane="6" heatid="22002" points="273" />
                <RESULT resultid="576" eventid="28" swimtime="00:00:31.93" lane="5" heatid="28003" points="339" />
                <RESULT resultid="577" eventid="40" swimtime="00:00:31.61" lane="8" heatid="40002" points="289" />
                <RESULT resultid="578" eventid="44" swimtime="00:00:41.92" lane="5" heatid="44001" points="237" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124" birthdate="2011-01-01" gender="M" lastname="Fabian" firstname="Constantin" license="430675" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:05.73" heatid="2005" lane="7" />
                <ENTRY eventid="12" entrytime="00:01:00.30" heatid="12004" lane="8" />
                <ENTRY eventid="24" entrytime="00:02:28.88" heatid="24003" lane="2" />
                <ENTRY eventid="38" entrytime="00:02:38.32" heatid="38001" lane="5" />
                <ENTRY eventid="46" entrytime="00:05:49.99" heatid="46001" lane="3" />
                <ENTRY eventid="15" entrytime="00:01:05.22" heatid="15001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="579" eventid="2" swimtime="00:01:05.22" lane="7" heatid="2005" points="435" />
                <RESULT resultid="580" eventid="12" swimtime="00:01:00.31" lane="8" heatid="12004" points="455" />
                <RESULT resultid="822" eventid="15" swimtime="00:01:05.39" lane="2" heatid="15001" points="432" />
                <RESULT resultid="581" eventid="24" swimtime="00:02:33.73" lane="2" heatid="24003" points="407">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="582" eventid="38" swimtime="00:02:31.50" lane="5" heatid="38001" points="386">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="583" eventid="46" swimtime="00:04:39.56" lane="3" heatid="46001" points="487">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.76" />
                    <SPLIT distance="200" swimtime="00:02:18.37" />
                    <SPLIT distance="300" swimtime="00:03:29.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125" birthdate="2012-01-01" gender="F" lastname="Kotelnytska" firstname="Daria" license="455829" nation="UKR">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:14.93" heatid="1002" lane="8" />
                <ENTRY eventid="7" entrytime="00:02:54.44" heatid="7001" lane="3" />
                <ENTRY eventid="23" entrytime="00:02:37.80" heatid="23004" lane="8" />
                <ENTRY eventid="27" entrytime="00:00:37.23" heatid="27002" lane="2" />
                <ENTRY eventid="37" entrytime="00:03:11.49" heatid="37001" lane="5" />
                <ENTRY eventid="45" entrytime="00:05:14.44" heatid="45002" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="584" eventid="1" swimtime="00:01:14.43" lane="8" heatid="1002" points="407" />
                <RESULT resultid="585" eventid="7" swimtime="00:02:39.37" lane="3" heatid="7001" points="461">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="586" eventid="23" swimtime="00:02:38.86" lane="8" heatid="23004" points="500">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="587" eventid="27" swimtime="00:00:33.56" lane="2" heatid="27002" points="385" />
                <RESULT resultid="588" eventid="37" swimtime="00:02:54.32" lane="5" heatid="37001" points="341">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="589" eventid="45" swimtime="00:04:59.74" lane="5" heatid="45002" points="484">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="200" swimtime="00:02:28.49" />
                    <SPLIT distance="300" swimtime="00:03:45.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="126" birthdate="2013-01-01" gender="M" lastname="Lüddecke" firstname="Emil" license="463238" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:44.41" heatid="2001" lane="3" />
                <ENTRY eventid="6" entrytime="00:02:05.66" heatid="6003" lane="1" />
                <ENTRY eventid="26" entrytime="00:00:00.00" heatid="26002" lane="7" />
                <ENTRY eventid="36" entrytime="00:01:19.24" heatid="36003" lane="8" />
                <ENTRY eventid="42" entrytime="00:00:00.00" heatid="42001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="590" eventid="2" swimtime="00:01:30.68" lane="3" heatid="2001" points="162" />
                <RESULT resultid="591" eventid="6" swimtime="00:01:40.00" lane="1" heatid="6003" points="184" />
                <RESULT resultid="592" eventid="26" swimtime="00:21:21.30" lane="7" heatid="26002" points="313">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.91" />
                    <SPLIT distance="200" swimtime="00:02:42.86" />
                    <SPLIT distance="300" swimtime="00:04:08.86" />
                    <SPLIT distance="400" swimtime="00:05:34.80" />
                    <SPLIT distance="500" swimtime="00:07:00.66" />
                    <SPLIT distance="600" swimtime="00:08:26.58" />
                    <SPLIT distance="700" swimtime="00:09:52.53" />
                    <SPLIT distance="800" swimtime="00:11:19.43" />
                    <SPLIT distance="900" swimtime="00:12:46.72" />
                    <SPLIT distance="1000" swimtime="00:14:13.76" />
                    <SPLIT distance="1100" swimtime="00:15:39.53" />
                    <SPLIT distance="1200" swimtime="00:17:06.44" />
                    <SPLIT distance="1300" swimtime="00:18:32.21" />
                    <SPLIT distance="1400" swimtime="00:19:58.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="593" eventid="36" swimtime="00:01:19.58" lane="8" heatid="36003" points="272" />
                <RESULT resultid="594" eventid="42" swimtime="00:06:23.45" lane="4" heatid="42001" points="252">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.90" />
                    <SPLIT distance="200" swimtime="00:03:11.17" />
                    <SPLIT distance="300" swimtime="00:05:02.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="127" birthdate="2012-01-01" gender="F" lastname="Vogt" firstname="Hilleda Sigune" license="442521" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:29.37" heatid="5002" lane="2" />
                <ENTRY eventid="11" entrytime="00:01:11.98" heatid="11002" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:56.01" heatid="23001" lane="6" />
                <ENTRY eventid="35" entrytime="00:01:24.45" heatid="35002" lane="1" />
                <ENTRY eventid="45" entrytime="00:05:28.10" heatid="45002" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="595" eventid="5" swimtime="00:01:30.72" lane="2" heatid="5002" points="353" />
                <RESULT resultid="596" eventid="11" swimtime="00:01:12.34" lane="5" heatid="11002" points="365" />
                <RESULT resultid="597" eventid="23" swimtime="00:02:53.14" lane="6" heatid="23001" points="386">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="598" eventid="35" swimtime="00:01:21.05" lane="1" heatid="35002" points="350" />
                <RESULT resultid="599" eventid="45" swimtime="00:05:26.52" lane="6" heatid="45002" points="374">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.40" />
                    <SPLIT distance="200" swimtime="00:02:39.88" />
                    <SPLIT distance="300" swimtime="00:04:04.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128" birthdate="2007-01-01" gender="F" lastname="Koch" firstname="Jette" license="369289" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:11.85" heatid="5002" lane="4" />
                <ENTRY eventid="23" entrytime="00:02:25.88" heatid="23005" lane="6" />
                <ENTRY eventid="27" entrytime="00:00:30.42" heatid="27004" lane="4" />
                <ENTRY eventid="39" entrytime="00:00:28.59" heatid="39003" lane="5" />
                <ENTRY eventid="43" entrytime="00:00:33.57" heatid="43003" lane="5" />
                <ENTRY eventid="18" entrytime="00:01:14.94" heatid="18001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="600" eventid="5" swimtime="00:01:14.94" lane="4" heatid="5002" points="626" />
                <RESULT resultid="842" eventid="18" swimtime="00:01:14.56" lane="5" heatid="18001" points="636" />
                <RESULT resultid="601" eventid="23" swimtime="00:02:34.47" lane="6" heatid="23005" points="544">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="602" eventid="27" swimtime="00:00:31.52" lane="4" heatid="27004" points="465" />
                <RESULT resultid="603" eventid="39" swimtime="00:00:29.28" lane="5" heatid="39003" points="524" />
                <RESULT resultid="604" eventid="43" swimtime="00:00:34.44" lane="5" heatid="43003" points="606" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129" birthdate="2006-01-01" gender="F" lastname="Barth" firstname="Julia" license="329294" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:02.58" heatid="3003" lane="4" />
                <ENTRY eventid="9" entrytime="00:08:54.03" heatid="9000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="605" eventid="3" status="WDR" swimtime="00:00:00.00" lane="4" heatid="3003" />
                <RESULT resultid="606" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130" birthdate="2012-01-01" gender="F" lastname="Slach" firstname="Katharina" license="436752" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:15.36" heatid="1001" lane="4" />
                <ENTRY eventid="9" entrytime="00:10:22.22" heatid="9002" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:34.52" heatid="27002" lane="3" />
                <ENTRY eventid="39" entrytime="00:00:30.19" heatid="39002" lane="6" />
                <ENTRY eventid="45" entrytime="00:05:03.91" heatid="45003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="607" eventid="1" swimtime="00:01:17.44" lane="4" heatid="1001" points="361" />
                <RESULT resultid="608" eventid="9" swimtime="00:10:20.19" lane="2" heatid="9002" points="477">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.14" />
                    <SPLIT distance="200" swimtime="00:02:29.72" />
                    <SPLIT distance="300" swimtime="00:03:47.42" />
                    <SPLIT distance="400" swimtime="00:05:06.52" />
                    <SPLIT distance="500" swimtime="00:06:25.07" />
                    <SPLIT distance="600" swimtime="00:07:43.90" />
                    <SPLIT distance="700" swimtime="00:09:02.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="609" eventid="27" swimtime="00:00:33.62" lane="3" heatid="27002" points="383" />
                <RESULT resultid="610" eventid="39" swimtime="00:00:30.77" lane="6" heatid="39002" points="451" />
                <RESULT resultid="611" eventid="45" swimtime="00:04:58.74" lane="1" heatid="45003" points="489">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="200" swimtime="00:02:28.98" />
                    <SPLIT distance="300" swimtime="00:03:45.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="131" birthdate="2013-01-01" gender="F" lastname="Staack" firstname="Kiki Marlen" license="459682" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:35.56" heatid="1001" lane="1" />
                <ENTRY eventid="9" entrytime="00:00:00.00" heatid="9001" lane="3" />
                <ENTRY eventid="23" entrytime="00:02:57.28" heatid="23001" lane="7" />
                <ENTRY eventid="29" entrytime="00:03:40.00" heatid="29001" lane="2" />
                <ENTRY eventid="35" entrytime="00:01:38.50" heatid="35001" lane="2" />
                <ENTRY eventid="41" entrytime="00:00:00.00" heatid="41001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="612" eventid="1" swimtime="00:01:22.29" lane="1" heatid="1001" points="301" />
                <RESULT resultid="613" eventid="9" swimtime="00:10:53.86" lane="3" heatid="9001" points="407">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.09" />
                    <SPLIT distance="200" swimtime="00:02:35.11" />
                    <SPLIT distance="300" swimtime="00:03:58.06" />
                    <SPLIT distance="400" swimtime="00:05:21.81" />
                    <SPLIT distance="500" swimtime="00:06:46.61" />
                    <SPLIT distance="600" swimtime="00:08:12.64" />
                    <SPLIT distance="700" swimtime="00:09:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="614" eventid="23" swimtime="00:02:54.27" lane="7" heatid="23001" points="379">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="615" eventid="29" swimtime="00:03:22.41" lane="2" heatid="29001" points="313">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="616" eventid="35" swimtime="00:01:23.02" lane="2" heatid="35001" points="325" />
                <RESULT resultid="617" eventid="41" swimtime="00:06:14.82" lane="6" heatid="41001" points="350">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.09" />
                    <SPLIT distance="200" swimtime="00:03:07.57" />
                    <SPLIT distance="300" swimtime="00:04:54.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="132" birthdate="2012-01-01" gender="F" lastname="Gutiérrez Müller" firstname="Laia" license="476631" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:10.33" heatid="1004" lane="2" />
                <ENTRY eventid="9" entrytime="00:10:16.66" heatid="9002" lane="6" />
                <ENTRY eventid="23" entrytime="00:02:34.70" heatid="23004" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:31.55" heatid="27003" lane="4" />
                <ENTRY eventid="39" entrytime="00:00:30.16" heatid="39002" lane="3" />
                <ENTRY eventid="45" entrytime="00:04:51.78" heatid="45003" lane="3" />
                <ENTRY eventid="13" entrytime="00:01:09.13" heatid="13001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="618" eventid="1" swimtime="00:01:09.13" lane="2" heatid="1004" points="508" />
                <RESULT resultid="619" eventid="9" swimtime="00:10:06.59" lane="6" heatid="9002" points="510">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.56" />
                    <SPLIT distance="200" swimtime="00:02:27.94" />
                    <SPLIT distance="300" swimtime="00:03:44.40" />
                    <SPLIT distance="400" swimtime="00:05:01.70" />
                    <SPLIT distance="500" swimtime="00:06:18.87" />
                    <SPLIT distance="600" swimtime="00:07:36.00" />
                    <SPLIT distance="700" swimtime="00:08:52.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="805" eventid="13" swimtime="00:01:09.16" lane="3" heatid="13001" points="507" />
                <RESULT resultid="620" eventid="23" swimtime="00:02:39.46" lane="2" heatid="23004" points="494">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="621" eventid="27" swimtime="00:00:30.90" lane="4" heatid="27003" points="494" />
                <RESULT resultid="622" eventid="39" swimtime="00:00:29.76" lane="3" heatid="39002" points="499" />
                <RESULT resultid="623" eventid="45" swimtime="00:04:55.88" lane="3" heatid="45003" points="503">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.97" />
                    <SPLIT distance="200" swimtime="00:02:24.66" />
                    <SPLIT distance="300" swimtime="00:03:41.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="133" birthdate="2005-01-01" gender="F" lastname="Braun" firstname="Lara" license="384947" nation="GER">
              <ENTRIES>
                <ENTRY eventid="25" entrytime="00:17:02.36" heatid="25000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="624" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="134" birthdate="2012-01-01" gender="F" lastname="Mühlbauer" firstname="Laura Charlotte" license="449363" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:22.81" heatid="1001" lane="6" />
                <ENTRY eventid="7" entrytime="00:02:39.18" heatid="7002" lane="8" />
                <ENTRY eventid="23" entrytime="00:02:46.63" heatid="23002" lane="2" />
                <ENTRY eventid="35" entrytime="00:01:12.03" heatid="35003" lane="2" />
                <ENTRY eventid="41" entrytime="00:05:56.65" heatid="41002" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="625" eventid="1" swimtime="00:01:18.81" lane="6" heatid="1001" points="343" />
                <RESULT resultid="626" eventid="7" swimtime="00:02:39.09" lane="8" heatid="7002" points="463">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="627" eventid="23" swimtime="00:02:41.42" lane="2" heatid="23002" points="476">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="628" eventid="35" swimtime="00:01:13.71" lane="2" heatid="35003" points="465" />
                <RESULT resultid="629" eventid="41" swimtime="00:05:50.05" lane="7" heatid="41002" points="430">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.44" />
                    <SPLIT distance="200" swimtime="00:02:51.45" />
                    <SPLIT distance="300" swimtime="00:04:31.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="135" birthdate="2009-01-01" gender="M" lastname="Tunc" firstname="Leander-Tharus" license="398946" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:03.00" heatid="2004" lane="3" />
                <ENTRY eventid="10" entrytime="00:09:41.98" heatid="10002" lane="7" />
                <ENTRY eventid="40" entrytime="00:00:26.95" heatid="40004" lane="7" />
                <ENTRY eventid="44" entrytime="00:00:33.93" heatid="44003" lane="8" />
                <ENTRY eventid="16" entrytime="00:01:02.08" heatid="16001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="630" eventid="2" swimtime="00:01:02.08" lane="3" heatid="2004" points="505" />
                <RESULT resultid="631" eventid="10" swimtime="00:10:00.60" lane="7" heatid="10002" points="426">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="200" swimtime="00:02:23.17" />
                    <SPLIT distance="300" swimtime="00:03:38.76" />
                    <SPLIT distance="400" swimtime="00:04:55.82" />
                    <SPLIT distance="500" swimtime="00:06:13.29" />
                    <SPLIT distance="600" swimtime="00:07:31.53" />
                    <SPLIT distance="700" swimtime="00:08:48.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="831" eventid="16" swimtime="00:01:01.97" lane="7" heatid="16001" points="508" />
                <RESULT resultid="632" eventid="40" swimtime="00:00:26.97" lane="7" heatid="40004" points="466" />
                <RESULT resultid="633" eventid="44" swimtime="00:00:33.48" lane="8" heatid="44003" points="465" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="136" birthdate="2010-01-01" gender="F" lastname="Werner" firstname="Lilli" license="430319" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:20.71" heatid="3002" lane="7" />
                <ENTRY eventid="23" entrytime="00:02:37.93" heatid="23003" lane="4" />
                <ENTRY eventid="29" entrytime="00:02:48.93" heatid="29002" lane="6" />
                <ENTRY eventid="35" entrytime="00:01:12.59" heatid="35005" lane="7" />
                <ENTRY eventid="41" entrytime="00:05:48.72" heatid="41002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="634" eventid="3" swimtime="00:02:31.95" lane="7" heatid="3002" points="402">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="635" eventid="23" swimtime="00:02:45.03" lane="4" heatid="23003" points="446">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="636" eventid="29" swimtime="00:03:05.83" lane="6" heatid="29002" points="405">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="637" eventid="35" swimtime="00:01:19.40" lane="7" heatid="35005" points="372" />
                <RESULT resultid="638" eventid="41" swimtime="00:05:54.09" lane="2" heatid="41002" points="416">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.16" />
                    <SPLIT distance="200" swimtime="00:02:55.11" />
                    <SPLIT distance="300" swimtime="00:04:33.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="137" birthdate="2010-01-01" gender="F" lastname="Barth" firstname="Lisa" license="377094" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:04.63" heatid="1002" lane="5" />
                <ENTRY eventid="9" entrytime="00:09:25.53" heatid="9000" lane="0" />
                <ENTRY eventid="27" entrytime="00:00:29.66" heatid="27005" lane="1" />
                <ENTRY eventid="35" entrytime="00:01:09.19" heatid="35004" lane="3" />
                <ENTRY eventid="39" entrytime="00:00:29.48" heatid="39003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="639" eventid="1" status="WDR" swimtime="00:00:00.00" lane="5" heatid="1002" />
                <RESULT resultid="640" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
                <RESULT resultid="641" eventid="27" status="WDR" swimtime="00:00:00.00" lane="1" heatid="27005" />
                <RESULT resultid="642" eventid="35" status="WDR" swimtime="00:00:00.00" lane="3" heatid="35004" />
                <RESULT resultid="643" eventid="39" status="WDR" swimtime="00:00:00.00" lane="1" heatid="39003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="138" birthdate="2010-01-01" gender="F" lastname="Adam" firstname="Lotta" license="414440" nation="GER">
              <ENTRIES>
                <ENTRY eventid="9" entrytime="00:09:15.05" heatid="9002" lane="5" />
                <ENTRY eventid="25" entrytime="00:17:44.57" heatid="25001" lane="4" />
                <ENTRY eventid="35" entrytime="00:01:08.57" heatid="35003" lane="5" />
                <ENTRY eventid="41" entrytime="00:05:14.06" heatid="41002" lane="5" />
                <ENTRY eventid="47" entrytime="00:01:11.30" heatid="47001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="644" eventid="9" swimtime="00:09:21.57" lane="5" heatid="9002" points="643">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                    <SPLIT distance="200" swimtime="00:02:15.47" />
                    <SPLIT distance="300" swimtime="00:03:25.55" />
                    <SPLIT distance="400" swimtime="00:04:36.11" />
                    <SPLIT distance="500" swimtime="00:05:47.05" />
                    <SPLIT distance="600" swimtime="00:06:58.62" />
                    <SPLIT distance="700" swimtime="00:08:10.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="645" eventid="25" swimtime="00:18:05.06" lane="4" heatid="25001" points="610">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.59" />
                    <SPLIT distance="200" swimtime="00:02:19.11" />
                    <SPLIT distance="300" swimtime="00:03:30.17" />
                    <SPLIT distance="400" swimtime="00:04:41.00" />
                    <SPLIT distance="500" swimtime="00:05:52.38" />
                    <SPLIT distance="600" swimtime="00:07:05.22" />
                    <SPLIT distance="700" swimtime="00:08:18.56" />
                    <SPLIT distance="800" swimtime="00:09:31.38" />
                    <SPLIT distance="900" swimtime="00:10:45.08" />
                    <SPLIT distance="1000" swimtime="00:11:58.53" />
                    <SPLIT distance="1100" swimtime="00:13:11.98" />
                    <SPLIT distance="1200" swimtime="00:14:25.50" />
                    <SPLIT distance="1300" swimtime="00:15:39.57" />
                    <SPLIT distance="1400" swimtime="00:16:53.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="646" eventid="35" swimtime="00:01:11.30" lane="5" heatid="35003" points="514" />
                <RESULT resultid="647" eventid="41" swimtime="00:05:20.59" lane="5" heatid="41002" points="560">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.91" />
                    <SPLIT distance="200" swimtime="00:02:40.85" />
                    <SPLIT distance="300" swimtime="00:04:09.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="892" eventid="47" swimtime="00:01:11.42" lane="2" heatid="47001" points="511" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="139" birthdate="2005-01-01" gender="M" lastname="Schöttge" firstname="Luca" license="324418" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:00:57.68" heatid="2005" lane="5" />
                <ENTRY eventid="8" entrytime="00:02:04.51" heatid="8003" lane="5" />
                <ENTRY eventid="24" entrytime="00:02:04.44" heatid="24000" lane="0" />
                <ENTRY eventid="36" entrytime="00:00:57.86" heatid="36002" lane="4" />
                <ENTRY eventid="38" entrytime="00:02:06.36" heatid="38002" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="648" eventid="2" status="WDR" swimtime="00:00:00.00" lane="5" heatid="2005" />
                <RESULT resultid="649" eventid="8" status="WDR" swimtime="00:00:00.00" lane="5" heatid="8003" />
                <RESULT resultid="650" eventid="24" status="WDR" swimtime="00:00:00.00" lane="0" heatid="24000" />
                <RESULT resultid="651" eventid="36" status="WDR" swimtime="00:00:00.00" lane="4" heatid="36002" />
                <RESULT resultid="652" eventid="38" status="WDR" swimtime="00:00:00.00" lane="6" heatid="38002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140" birthdate="2013-01-01" gender="F" lastname="Preuß" firstname="Marie" license="442524" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:24.51" heatid="1001" lane="2" />
                <ENTRY eventid="9" entrytime="00:00:00.00" heatid="9001" lane="4" />
                <ENTRY eventid="23" entrytime="00:02:50.75" heatid="23002" lane="1" />
                <ENTRY eventid="29" entrytime="00:03:15.84" heatid="29001" lane="4" />
                <ENTRY eventid="35" entrytime="00:01:37.02" heatid="35001" lane="6" />
                <ENTRY eventid="41" entrytime="00:00:00.00" heatid="41001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="653" eventid="1" swimtime="00:01:20.54" lane="2" heatid="1001" points="321" />
                <RESULT resultid="654" eventid="9" swimtime="00:11:15.85" lane="4" heatid="9001" points="369">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.50" />
                    <SPLIT distance="200" swimtime="00:02:45.28" />
                    <SPLIT distance="300" swimtime="00:04:11.84" />
                    <SPLIT distance="400" swimtime="00:05:37.98" />
                    <SPLIT distance="500" swimtime="00:07:05.28" />
                    <SPLIT distance="600" swimtime="00:08:31.31" />
                    <SPLIT distance="700" swimtime="00:09:56.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="655" eventid="23" swimtime="00:02:47.80" lane="1" heatid="23002" points="424">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="656" eventid="29" swimtime="00:03:12.43" lane="4" heatid="29001" points="365">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="657" eventid="35" swimtime="00:01:21.43" lane="6" heatid="35001" points="345" />
                <RESULT resultid="658" eventid="41" swimtime="00:05:55.78" lane="3" heatid="41001" points="410">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                    <SPLIT distance="200" swimtime="00:02:56.03" />
                    <SPLIT distance="300" swimtime="00:04:37.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="141" birthdate="2011-01-01" gender="F" lastname="Himmel" firstname="Marlene" license="442520" nation="GER">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:02:34.33" heatid="7002" lane="7" />
                <ENTRY eventid="11" entrytime="00:01:05.95" heatid="11004" lane="8" />
                <ENTRY eventid="23" entrytime="00:02:48.11" heatid="23002" lane="7" />
                <ENTRY eventid="35" entrytime="00:01:12.72" heatid="35004" lane="7" />
                <ENTRY eventid="45" entrytime="00:05:09.40" heatid="45002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="659" eventid="7" swimtime="00:02:36.15" lane="7" heatid="7002" points="490">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="660" eventid="11" swimtime="00:01:05.73" lane="8" heatid="11004" points="486" />
                <RESULT resultid="661" eventid="23" swimtime="00:02:44.25" lane="7" heatid="23002" points="452">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="662" eventid="35" swimtime="00:01:14.09" lane="7" heatid="35004" points="458" />
                <RESULT resultid="663" eventid="45" swimtime="00:05:06.69" lane="4" heatid="45002" points="452">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="200" swimtime="00:02:31.14" />
                    <SPLIT distance="300" swimtime="00:03:49.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="142" birthdate="2009-01-01" gender="M" lastname="Nebelung" firstname="Mattis" license="369734" nation="GER">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:02:17.82" heatid="8003" lane="8" />
                <ENTRY eventid="26" entrytime="00:17:55.79" heatid="26002" lane="5" />
                <ENTRY eventid="42" entrytime="00:05:09.19" heatid="42003" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="664" eventid="8" swimtime="00:02:24.42" lane="8" heatid="8003" points="465">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="665" eventid="26" swimtime="00:17:33.70" lane="5" heatid="26002" points="564">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.18" />
                    <SPLIT distance="200" swimtime="00:02:16.07" />
                    <SPLIT distance="300" swimtime="00:03:27.37" />
                    <SPLIT distance="400" swimtime="00:04:38.30" />
                    <SPLIT distance="500" swimtime="00:05:49.45" />
                    <SPLIT distance="600" swimtime="00:07:00.16" />
                    <SPLIT distance="700" swimtime="00:08:10.90" />
                    <SPLIT distance="800" swimtime="00:09:21.58" />
                    <SPLIT distance="900" swimtime="00:10:32.15" />
                    <SPLIT distance="1000" swimtime="00:11:43.09" />
                    <SPLIT distance="1100" swimtime="00:12:53.91" />
                    <SPLIT distance="1200" swimtime="00:14:05.17" />
                    <SPLIT distance="1300" swimtime="00:15:16.36" />
                    <SPLIT distance="1400" swimtime="00:16:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="666" eventid="42" swimtime="00:05:02.65" lane="5" heatid="42003" points="514">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="200" swimtime="00:02:24.61" />
                    <SPLIT distance="300" swimtime="00:03:56.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143" birthdate="2014-01-01" gender="M" lastname="Kraus" firstname="Maximilian" license="443519" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:30.80" heatid="2001" lane="4" />
                <ENTRY eventid="6" entrytime="00:01:45.46" heatid="6001" lane="7" />
                <ENTRY eventid="26" entrytime="00:00:00.00" heatid="26001" lane="4" />
                <ENTRY eventid="36" entrytime="00:01:19.44" heatid="36002" lane="8" />
                <ENTRY eventid="42" entrytime="00:00:00.00" heatid="42002" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="667" eventid="2" swimtime="00:01:21.00" lane="4" heatid="2001" points="227" />
                <RESULT resultid="668" eventid="6" swimtime="00:01:44.14" lane="7" heatid="6001" points="162" />
                <RESULT resultid="669" eventid="26" swimtime="00:19:54.10" lane="4" heatid="26001" points="387">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.88" />
                    <SPLIT distance="200" swimtime="00:02:32.62" />
                    <SPLIT distance="300" swimtime="00:03:52.10" />
                    <SPLIT distance="400" swimtime="00:05:12.07" />
                    <SPLIT distance="500" swimtime="00:06:32.68" />
                    <SPLIT distance="600" swimtime="00:07:53.49" />
                    <SPLIT distance="700" swimtime="00:09:13.37" />
                    <SPLIT distance="800" swimtime="00:10:33.08" />
                    <SPLIT distance="900" swimtime="00:11:53.65" />
                    <SPLIT distance="1000" swimtime="00:13:16.07" />
                    <SPLIT distance="1100" swimtime="00:14:37.18" />
                    <SPLIT distance="1200" swimtime="00:15:58.00" />
                    <SPLIT distance="1300" swimtime="00:17:18.33" />
                    <SPLIT distance="1400" swimtime="00:18:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="670" eventid="36" swimtime="00:01:21.87" lane="8" heatid="36002" points="250" />
                <RESULT resultid="671" eventid="42" swimtime="00:06:08.14" lane="7" heatid="42002" points="285">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="200" swimtime="00:02:59.85" />
                    <SPLIT distance="300" swimtime="00:04:50.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144" birthdate="2010-01-01" gender="M" lastname="Wiemer" firstname="Maximilian" license="409856" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:23.68" heatid="6003" lane="6" />
                <ENTRY eventid="12" entrytime="00:00:56.58" heatid="12004" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:27.79" heatid="28005" lane="4" />
                <ENTRY eventid="40" entrytime="00:00:26.74" heatid="40004" lane="3" />
                <ENTRY eventid="46" entrytime="00:04:27.79" heatid="46003" lane="7" />
                <ENTRY eventid="19" entrytime="00:01:16.55" heatid="19001" lane="7" />
                <ENTRY eventid="33" entrytime="00:00:57.55" heatid="33001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="672" eventid="6" swimtime="00:01:16.55" lane="6" heatid="6003" points="410" />
                <RESULT resultid="673" eventid="12" swimtime="00:00:57.55" lane="2" heatid="12004" points="524" />
                <RESULT resultid="850" eventid="19" swimtime="00:01:17.20" lane="7" heatid="19001" points="399" />
                <RESULT resultid="674" eventid="28" swimtime="00:00:28.15" lane="4" heatid="28005" points="495" />
                <RESULT resultid="872" eventid="33" swimtime="00:00:56.69" lane="5" heatid="33001" points="548" />
                <RESULT resultid="675" eventid="40" swimtime="00:00:26.68" lane="3" heatid="40004" points="481" />
                <RESULT resultid="676" eventid="46" swimtime="00:05:24.80" lane="7" heatid="46003" points="311">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="200" swimtime="00:02:34.90" />
                    <SPLIT distance="300" swimtime="00:04:02.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145" birthdate="2013-01-01" gender="M" lastname="Deckenbach" firstname="Paul" license="453535" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:28.54" heatid="2002" lane="7" />
                <ENTRY eventid="6" entrytime="00:01:28.65" heatid="6003" lane="2" />
                <ENTRY eventid="26" entrytime="00:00:00.00" heatid="26002" lane="1" />
                <ENTRY eventid="36" entrytime="00:01:21.61" heatid="36001" lane="6" />
                <ENTRY eventid="42" entrytime="00:00:00.00" heatid="42002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="677" eventid="2" swimtime="00:01:20.32" lane="7" heatid="2002" points="233" />
                <RESULT resultid="678" eventid="6" swimtime="00:01:26.79" lane="2" heatid="6003" points="281" />
                <RESULT resultid="679" eventid="26" swimtime="00:21:38.78" lane="1" heatid="26002" points="301">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="200" swimtime="00:02:42.69" />
                    <SPLIT distance="300" swimtime="00:04:10.55" />
                    <SPLIT distance="400" swimtime="00:05:36.81" />
                    <SPLIT distance="500" swimtime="00:07:03.92" />
                    <SPLIT distance="600" swimtime="00:08:31.09" />
                    <SPLIT distance="700" swimtime="00:09:58.16" />
                    <SPLIT distance="800" swimtime="00:11:25.96" />
                    <SPLIT distance="900" swimtime="00:12:53.38" />
                    <SPLIT distance="1000" swimtime="00:14:20.84" />
                    <SPLIT distance="1100" swimtime="00:15:48.61" />
                    <SPLIT distance="1200" swimtime="00:17:17.67" />
                    <SPLIT distance="1300" swimtime="00:18:46.68" />
                    <SPLIT distance="1400" swimtime="00:20:14.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="680" eventid="36" swimtime="00:01:21.01" lane="6" heatid="36001" points="258" />
                <RESULT resultid="681" eventid="42" swimtime="00:05:59.58" lane="2" heatid="42002" points="306">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.23" />
                    <SPLIT distance="200" swimtime="00:02:58.35" />
                    <SPLIT distance="300" swimtime="00:04:35.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="146" birthdate="2010-01-01" gender="M" lastname="Schmidt" firstname="Paul" license="409854" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:07.21" heatid="2003" lane="7" />
                <ENTRY eventid="10" entrytime="00:09:50.55" heatid="10002" lane="8" />
                <ENTRY eventid="24" entrytime="00:02:26.31" heatid="24003" lane="5" />
                <ENTRY eventid="28" entrytime="00:00:00.00" heatid="28001" lane="3" />
                <ENTRY eventid="36" entrytime="00:01:12.22" heatid="36003" lane="7" />
                <ENTRY eventid="42" entrytime="00:05:12.78" heatid="42003" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="682" eventid="2" swimtime="00:01:06.67" lane="7" heatid="2003" points="408" />
                <RESULT resultid="683" eventid="10" swimtime="00:09:58.74" lane="8" heatid="10002" points="430">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="200" swimtime="00:02:24.66" />
                    <SPLIT distance="300" swimtime="00:03:39.55" />
                    <SPLIT distance="400" swimtime="00:04:54.96" />
                    <SPLIT distance="500" swimtime="00:06:11.79" />
                    <SPLIT distance="600" swimtime="00:07:28.80" />
                    <SPLIT distance="700" swimtime="00:08:45.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="684" eventid="24" swimtime="00:02:28.44" lane="5" heatid="24003" points="452">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="685" eventid="28" swimtime="00:00:29.41" lane="3" heatid="28001" points="434" />
                <RESULT resultid="686" eventid="36" swimtime="00:01:14.26" lane="7" heatid="36003" points="335" />
                <RESULT resultid="687" eventid="42" swimtime="00:05:22.56" lane="3" heatid="42003" points="424">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.22" />
                    <SPLIT distance="200" swimtime="00:02:37.54" />
                    <SPLIT distance="300" swimtime="00:04:08.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147" birthdate="2014-01-01" gender="F" lastname="Himmel" firstname="Paula" license="453672" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:22.23" heatid="1001" lane="3" />
                <ENTRY eventid="9" entrytime="00:00:00.00" heatid="9001" lane="6" />
                <ENTRY eventid="23" entrytime="00:02:57.01" heatid="23001" lane="2" />
                <ENTRY eventid="29" entrytime="00:03:40.00" heatid="29001" lane="6" />
                <ENTRY eventid="35" entrytime="00:01:33.74" heatid="35001" lane="5" />
                <ENTRY eventid="41" entrytime="00:00:00.00" heatid="41001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="688" eventid="1" swimtime="00:01:24.51" lane="3" heatid="1001" points="278" />
                <RESULT resultid="689" eventid="9" swimtime="00:11:22.89" lane="6" heatid="9001" points="357">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="200" swimtime="00:02:46.21" />
                    <SPLIT distance="300" swimtime="00:04:13.61" />
                    <SPLIT distance="400" swimtime="00:05:40.69" />
                    <SPLIT distance="500" swimtime="00:07:06.90" />
                    <SPLIT distance="600" swimtime="00:08:33.33" />
                    <SPLIT distance="700" swimtime="00:09:59.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="690" eventid="23" swimtime="00:02:59.61" lane="2" heatid="23001" points="346">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="691" eventid="29" swimtime="00:03:37.06" lane="6" heatid="29001" points="254">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="692" eventid="35" swimtime="00:01:23.69" lane="5" heatid="35001" points="318" />
                <RESULT resultid="693" eventid="41" swimtime="00:06:23.08" lane="5" heatid="41001" points="328">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.03" />
                    <SPLIT distance="200" swimtime="00:03:07.14" />
                    <SPLIT distance="300" swimtime="00:05:01.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="148" birthdate="2009-01-01" gender="F" lastname="Fertig" firstname="Pauline" license="370140" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:16.58" heatid="3002" lane="5" />
                <ENTRY eventid="9" entrytime="00:10:44.40" heatid="9002" lane="7" />
                <ENTRY eventid="41" entrytime="00:05:45.33" heatid="41002" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="694" eventid="3" swimtime="00:02:15.50" lane="5" heatid="3002" points="568">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="695" eventid="9" swimtime="00:10:03.94" lane="7" heatid="9002" points="517">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="200" swimtime="00:02:26.30" />
                    <SPLIT distance="300" swimtime="00:03:42.59" />
                    <SPLIT distance="400" swimtime="00:05:01.00" />
                    <SPLIT distance="500" swimtime="00:06:17.90" />
                    <SPLIT distance="600" swimtime="00:07:35.52" />
                    <SPLIT distance="700" swimtime="00:08:50.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="696" eventid="41" swimtime="00:05:35.23" lane="6" heatid="41002" points="490">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="200" swimtime="00:02:38.03" />
                    <SPLIT distance="300" swimtime="00:04:20.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149" birthdate="2008-01-01" gender="M" lastname="Bordas" firstname="Roland" license="388751" nation="GER">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:02:15.87" heatid="8003" lane="7" />
                <ENTRY eventid="12" entrytime="00:00:54.22" heatid="12005" lane="5" />
                <ENTRY eventid="24" entrytime="00:02:13.17" heatid="24004" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:26.44" heatid="28006" lane="2" />
                <ENTRY eventid="34" entrytime="00:00:54.92" heatid="34001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="697" eventid="8" swimtime="00:02:13.67" lane="7" heatid="8003" points="586">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="698" eventid="12" swimtime="00:00:54.92" lane="5" heatid="12005" points="603" />
                <RESULT resultid="699" eventid="24" swimtime="00:02:13.62" lane="3" heatid="24004" points="621">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="700" eventid="28" swimtime="00:00:27.29" lane="2" heatid="28006" points="543" />
                <RESULT resultid="884" eventid="34" swimtime="00:00:55.07" lane="2" heatid="34001" points="598" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150" birthdate="2006-01-01" gender="F" lastname="Schlump" firstname="Seike" license="346179" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:01.83" heatid="1003" lane="4" />
                <ENTRY eventid="3" entrytime="00:02:04.42" heatid="3003" lane="3" />
                <ENTRY eventid="37" entrytime="00:02:15.91" heatid="37002" lane="5" />
                <ENTRY eventid="14" entrytime="00:01:04.10" heatid="14000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="701" eventid="1" swimtime="00:01:04.10" lane="4" heatid="1003" points="637" />
                <RESULT resultid="702" eventid="3" swimtime="00:02:14.67" lane="3" heatid="3003" points="578">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="812" eventid="14" status="WDR" swimtime="00:00:00.00" lane="0" heatid="14000" />
                <RESULT resultid="703" eventid="37" swimtime="00:02:20.90" lane="5" heatid="37002" points="646">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="151" birthdate="2014-01-01" gender="F" lastname="Franke" firstname="Selina" license="449356" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:41.12" heatid="1001" lane="8" />
                <ENTRY eventid="9" entrytime="00:00:00.00" heatid="9001" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:53.11" heatid="23001" lane="5" />
                <ENTRY eventid="29" entrytime="00:03:30.00" heatid="29001" lane="3" />
                <ENTRY eventid="35" entrytime="00:01:18.11" heatid="35002" lane="3" />
                <ENTRY eventid="41" entrytime="00:00:00.00" heatid="41001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="704" eventid="1" swimtime="00:01:31.95" lane="8" heatid="1001" points="216" />
                <RESULT resultid="705" eventid="9" swimtime="00:11:19.02" lane="5" heatid="9001" points="363">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="200" swimtime="00:02:43.09" />
                    <SPLIT distance="300" swimtime="00:04:10.20" />
                    <SPLIT distance="400" swimtime="00:05:37.50" />
                    <SPLIT distance="500" swimtime="00:07:05.48" />
                    <SPLIT distance="600" swimtime="00:08:32.01" />
                    <SPLIT distance="700" swimtime="00:09:57.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="706" eventid="23" swimtime="00:02:52.07" lane="5" heatid="23001" points="393">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="707" eventid="29" swimtime="00:03:25.06" lane="3" heatid="29001" points="301">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="708" eventid="35" swimtime="00:01:17.91" lane="3" heatid="35002" points="394" />
                <RESULT resultid="709" eventid="41" swimtime="00:06:14.64" lane="2" heatid="41001" points="351">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.94" />
                    <SPLIT distance="200" swimtime="00:03:05.43" />
                    <SPLIT distance="300" swimtime="00:04:56.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="152" birthdate="2014-01-01" gender="F" lastname="Raguschke" firstname="Stella Shirly" license="469355" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:54.06" heatid="5001" lane="7" />
                <ENTRY eventid="11" entrytime="00:01:28.96" heatid="11001" lane="3" />
                <ENTRY eventid="21" entrytime="00:00:41.55" heatid="21001" lane="3" />
                <ENTRY eventid="27" entrytime="00:00:41.31" heatid="27001" lane="5" />
                <ENTRY eventid="39" entrytime="00:00:37.49" heatid="39001" lane="3" />
                <ENTRY eventid="43" entrytime="00:00:52.44" heatid="43001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="710" eventid="5" swimtime="00:01:41.18" lane="7" heatid="5001" points="254" />
                <RESULT resultid="711" eventid="11" swimtime="00:01:20.25" lane="3" heatid="11001" points="267" />
                <RESULT resultid="712" eventid="21" swimtime="00:00:41.46" lane="3" heatid="21001" points="271" />
                <RESULT resultid="713" eventid="27" swimtime="00:00:37.79" lane="5" heatid="27001" points="270" />
                <RESULT resultid="714" eventid="39" swimtime="00:00:36.77" lane="3" heatid="39001" points="264" />
                <RESULT resultid="715" eventid="43" swimtime="00:00:47.55" lane="3" heatid="43001" points="230" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="153" birthdate="2012-01-01" gender="F" lastname="Horn" firstname="Tessa" license="440188" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:19.31" heatid="3002" lane="6" />
                <ENTRY eventid="11" entrytime="00:01:04.40" heatid="11004" lane="1" />
                <ENTRY eventid="25" entrytime="00:19:52.46" heatid="25001" lane="3" />
                <ENTRY eventid="35" entrytime="00:01:15.64" heatid="35004" lane="8" />
                <ENTRY eventid="45" entrytime="00:04:52.32" heatid="45003" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="716" eventid="3" swimtime="00:02:18.99" lane="6" heatid="3002" points="526">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="717" eventid="11" swimtime="00:01:04.60" lane="1" heatid="11004" points="512" />
                <RESULT resultid="718" eventid="25" swimtime="00:19:01.54" lane="3" heatid="25001" points="524">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.30" />
                    <SPLIT distance="200" swimtime="00:02:26.61" />
                    <SPLIT distance="300" swimtime="00:03:42.37" />
                    <SPLIT distance="400" swimtime="00:04:58.67" />
                    <SPLIT distance="500" swimtime="00:06:15.38" />
                    <SPLIT distance="600" swimtime="00:07:31.82" />
                    <SPLIT distance="700" swimtime="00:08:48.83" />
                    <SPLIT distance="800" swimtime="00:10:05.70" />
                    <SPLIT distance="900" swimtime="00:11:22.00" />
                    <SPLIT distance="1000" swimtime="00:12:38.75" />
                    <SPLIT distance="1100" swimtime="00:13:55.19" />
                    <SPLIT distance="1200" swimtime="00:15:12.25" />
                    <SPLIT distance="1300" swimtime="00:16:29.35" />
                    <SPLIT distance="1400" swimtime="00:17:47.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="719" eventid="35" swimtime="00:01:15.38" lane="8" heatid="35004" points="435" />
                <RESULT resultid="720" eventid="45" swimtime="00:04:51.63" lane="6" heatid="45003" points="525">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.91" />
                    <SPLIT distance="200" swimtime="00:02:22.46" />
                    <SPLIT distance="300" swimtime="00:03:37.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154" birthdate="2013-01-01" gender="M" lastname="Schreiber" firstname="Toni" license="442728" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:30.00" heatid="2002" lane="1" />
                <ENTRY eventid="6" entrytime="00:01:40.48" heatid="6002" lane="7" />
                <ENTRY eventid="26" entrytime="00:00:00.00" heatid="26001" lane="5" />
                <ENTRY eventid="36" entrytime="00:01:14.76" heatid="36004" lane="1" />
                <ENTRY eventid="42" entrytime="00:00:00.00" heatid="42001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="721" eventid="2" swimtime="00:01:23.99" lane="1" heatid="2002" points="204" />
                <RESULT resultid="722" eventid="6" swimtime="00:01:38.77" lane="7" heatid="6002" points="190" />
                <RESULT resultid="723" eventid="26" swimtime="00:21:23.44" lane="5" heatid="26001" points="312">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.17" />
                    <SPLIT distance="200" swimtime="00:02:45.64" />
                    <SPLIT distance="300" swimtime="00:04:11.96" />
                    <SPLIT distance="400" swimtime="00:05:39.91" />
                    <SPLIT distance="500" swimtime="00:07:08.86" />
                    <SPLIT distance="600" swimtime="00:08:35.18" />
                    <SPLIT distance="700" swimtime="00:10:03.42" />
                    <SPLIT distance="800" swimtime="00:11:29.88" />
                    <SPLIT distance="900" swimtime="00:12:54.88" />
                    <SPLIT distance="1000" swimtime="00:14:21.70" />
                    <SPLIT distance="1100" swimtime="00:15:48.03" />
                    <SPLIT distance="1200" swimtime="00:17:12.83" />
                    <SPLIT distance="1300" swimtime="00:18:38.30" />
                    <SPLIT distance="1400" swimtime="00:20:02.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="724" eventid="36" swimtime="00:01:14.70" lane="1" heatid="36004" points="329" />
                <RESULT resultid="725" eventid="42" swimtime="00:06:07.47" lane="5" heatid="42001" points="287">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.30" />
                    <SPLIT distance="200" swimtime="00:03:00.01" />
                    <SPLIT distance="300" swimtime="00:04:50.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="155" birthdate="2014-01-01" gender="M" lastname="Schwedler" firstname="Willi" license="445877" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:31.59" heatid="2001" lane="5" />
                <ENTRY eventid="6" entrytime="00:01:38.89" heatid="6003" lane="7" />
                <ENTRY eventid="26" entrytime="00:00:00.00" heatid="26001" lane="3" />
                <ENTRY eventid="36" entrytime="00:01:20.72" heatid="36001" lane="4" />
                <ENTRY eventid="42" entrytime="00:00:00.00" heatid="42001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="726" eventid="2" swimtime="00:01:22.79" lane="5" heatid="2001" points="213" />
                <RESULT resultid="727" eventid="6" swimtime="00:01:37.10" lane="7" heatid="6003" points="201" />
                <RESULT resultid="728" eventid="26" swimtime="00:22:43.55" lane="3" heatid="26001" points="260">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.79" />
                    <SPLIT distance="200" swimtime="00:02:50.16" />
                    <SPLIT distance="300" swimtime="00:04:21.19" />
                    <SPLIT distance="400" swimtime="00:05:53.10" />
                    <SPLIT distance="500" swimtime="00:07:25.07" />
                    <SPLIT distance="600" swimtime="00:08:57.55" />
                    <SPLIT distance="700" swimtime="00:10:29.98" />
                    <SPLIT distance="800" swimtime="00:12:01.64" />
                    <SPLIT distance="900" swimtime="00:13:34.98" />
                    <SPLIT distance="1000" swimtime="00:15:07.90" />
                    <SPLIT distance="1100" swimtime="00:16:41.72" />
                    <SPLIT distance="1200" swimtime="00:18:13.63" />
                    <SPLIT distance="1300" swimtime="00:19:45.60" />
                    <SPLIT distance="1400" swimtime="00:21:16.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="729" eventid="36" swimtime="00:01:20.45" lane="4" heatid="36001" points="263" />
                <RESULT resultid="730" eventid="42" swimtime="00:06:11.66" lane="3" heatid="42001" points="277">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.59" />
                    <SPLIT distance="200" swimtime="00:03:03.42" />
                    <SPLIT distance="300" swimtime="00:04:48.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Riesa" nation="GER" region="12" code="3356">
          <ATHLETES>
            <ATHLETE athleteid="45" birthdate="2013-01-01" gender="M" lastname="Thomas" firstname="Florin" license="437788" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:21.00" heatid="2002" lane="6" />
                <ENTRY eventid="12" entrytime="00:01:08.02" heatid="12002" lane="7" />
                <ENTRY eventid="22" entrytime="00:00:37.93" heatid="22002" lane="8" />
                <ENTRY eventid="28" entrytime="00:00:35.01" heatid="28002" lane="4" />
                <ENTRY eventid="36" entrytime="00:01:22.37" heatid="36001" lane="2" />
                <ENTRY eventid="42" entrytime="00:05:53.09" heatid="42002" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="221" eventid="2" swimtime="00:01:17.14" lane="6" heatid="2002" points="263" />
                <RESULT resultid="222" eventid="12" swimtime="00:01:05.92" lane="7" heatid="12002" points="348" />
                <RESULT resultid="223" eventid="22" swimtime="00:00:37.22" lane="8" heatid="22002" points="253" />
                <RESULT resultid="224" eventid="28" swimtime="00:00:33.51" lane="4" heatid="28002" points="293" />
                <RESULT resultid="225" eventid="36" swimtime="00:01:20.01" lane="2" heatid="36001" points="268" />
                <RESULT resultid="226" eventid="42" swimtime="00:05:42.14" lane="4" heatid="42002" points="356">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.78" />
                    <SPLIT distance="200" swimtime="00:02:54.01" />
                    <SPLIT distance="300" swimtime="00:04:26.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="46" birthdate="2013-01-01" gender="M" lastname="Schäfer" firstname="Jonas" license="449096" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:34.07" heatid="4002" lane="2" />
                <ENTRY eventid="10" entrytime="00:11:27.72" heatid="10001" lane="8" />
                <ENTRY eventid="26" entrytime="00:21:32.08" heatid="26002" lane="2" />
                <ENTRY eventid="40" entrytime="00:00:31.88" heatid="40001" lane="4" />
                <ENTRY eventid="42" entrytime="00:06:14.77" heatid="42002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="227" eventid="4" swimtime="00:02:31.38" lane="2" heatid="4002" points="305">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="228" eventid="10" swimtime="00:10:41.94" lane="8" heatid="10001" points="349">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="200" swimtime="00:02:34.65" />
                    <SPLIT distance="300" swimtime="00:03:56.27" />
                    <SPLIT distance="400" swimtime="00:05:18.31" />
                    <SPLIT distance="500" swimtime="00:06:39.78" />
                    <SPLIT distance="600" swimtime="00:08:02.31" />
                    <SPLIT distance="700" swimtime="00:09:23.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="229" eventid="26" swimtime="00:20:29.07" lane="2" heatid="26002" points="355">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                    <SPLIT distance="200" swimtime="00:02:36.70" />
                    <SPLIT distance="300" swimtime="00:03:59.19" />
                    <SPLIT distance="400" swimtime="00:05:21.04" />
                    <SPLIT distance="500" swimtime="00:06:43.74" />
                    <SPLIT distance="600" swimtime="00:08:06.47" />
                    <SPLIT distance="700" swimtime="00:09:29.30" />
                    <SPLIT distance="800" swimtime="00:10:51.99" />
                    <SPLIT distance="900" swimtime="00:12:14.98" />
                    <SPLIT distance="1000" swimtime="00:13:36.79" />
                    <SPLIT distance="1100" swimtime="00:15:00.12" />
                    <SPLIT distance="1200" swimtime="00:16:23.08" />
                    <SPLIT distance="1300" swimtime="00:17:46.40" />
                    <SPLIT distance="1400" swimtime="00:19:09.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="230" eventid="40" swimtime="00:00:30.70" lane="4" heatid="40001" points="315" />
                <RESULT resultid="231" eventid="42" swimtime="00:06:02.49" lane="3" heatid="42002" points="299">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.25" />
                    <SPLIT distance="200" swimtime="00:03:01.47" />
                    <SPLIT distance="300" swimtime="00:04:46.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="47" birthdate="2013-01-01" gender="M" lastname="Mühlmann" firstname="Ole" license="446953" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:28.93" heatid="6002" lane="2" />
                <ENTRY eventid="12" entrytime="00:01:09.89" heatid="12001" lane="4" />
                <ENTRY eventid="22" entrytime="00:00:38.17" heatid="22001" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:34.97" heatid="28003" lane="8" />
                <ENTRY eventid="38" entrytime="00:03:56.83" heatid="38001" lane="7" />
                <ENTRY eventid="44" entrytime="00:00:40.40" heatid="44002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="232" eventid="6" swimtime="00:01:28.76" lane="2" heatid="6002" points="263" />
                <RESULT resultid="233" eventid="12" swimtime="00:01:09.76" lane="4" heatid="12001" points="294" />
                <RESULT resultid="234" eventid="22" swimtime="00:00:36.91" lane="4" heatid="22001" points="259" />
                <RESULT resultid="235" eventid="28" swimtime="00:00:33.51" lane="8" heatid="28003" points="293" />
                <RESULT resultid="236" eventid="38" status="DSQ" swimtime="00:03:12.96" lane="7" heatid="38001" comment="Der Sportler führte auf der Schwimmstrecke Wechselbeinbewegungen aus und schlug bei der 1. &amp; 3. Wende nicht mit beiden Händen gleichzeitig an.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="237" eventid="44" swimtime="00:00:39.85" lane="2" heatid="44002" points="276" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SSG Leipzig e.V." nation="GER" region="12" code="6466">
          <ATHLETES>
            <ATHLETE athleteid="13" birthdate="2006-01-01" gender="F" lastname="Schiffel" firstname="Aaliyah" license="348758" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:10.97" heatid="5003" lane="4" />
                <ENTRY eventid="23" entrytime="00:02:18.17" heatid="23005" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:29.39" heatid="27005" lane="2" />
                <ENTRY eventid="18" entrytime="00:01:11.87" heatid="18001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="54" eventid="5" swimtime="00:01:11.87" lane="4" heatid="5003" points="710" />
                <RESULT resultid="841" eventid="18" swimtime="00:01:11.72" lane="4" heatid="18001" points="714" />
                <RESULT resultid="55" eventid="23" swimtime="00:02:21.19" lane="4" heatid="23005" points="712">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="56" eventid="27" swimtime="00:00:29.18" lane="2" heatid="27005" points="586" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="14" birthdate="2010-01-01" gender="M" lastname="Belyavskiy" firstname="Alexander" license="426136" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:09:02.11" heatid="10002" lane="5" />
                <ENTRY eventid="24" entrytime="00:02:25.19" heatid="24003" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:28.38" heatid="28005" lane="3" />
                <ENTRY eventid="36" entrytime="00:01:07.80" heatid="36003" lane="6" />
                <ENTRY eventid="40" entrytime="00:00:27.24" heatid="40004" lane="1" />
                <ENTRY eventid="49" entrytime="00:01:07.71" heatid="49001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="57" eventid="10" swimtime="00:08:55.70" lane="5" heatid="10002" points="601">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.06" />
                    <SPLIT distance="200" swimtime="00:02:08.71" />
                    <SPLIT distance="300" swimtime="00:03:16.09" />
                    <SPLIT distance="400" swimtime="00:04:24.29" />
                    <SPLIT distance="500" swimtime="00:05:32.44" />
                    <SPLIT distance="600" swimtime="00:06:40.64" />
                    <SPLIT distance="700" swimtime="00:07:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="58" eventid="24" swimtime="00:02:23.03" lane="4" heatid="24003" points="506">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="59" eventid="28" swimtime="00:00:28.46" lane="3" heatid="28005" points="479" />
                <RESULT resultid="60" eventid="36" swimtime="00:01:07.71" lane="6" heatid="36003" points="442" />
                <RESULT resultid="61" eventid="40" swimtime="00:00:27.64" lane="1" heatid="40004" points="432" />
                <RESULT resultid="904" eventid="49" swimtime="00:01:06.38" lane="6" heatid="49001" points="469" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="15" birthdate="2011-01-01" gender="F" lastname="Hunger" firstname="Anna Franziska" license="428578" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:08.02" heatid="1003" lane="6" />
                <ENTRY eventid="5" entrytime="00:01:15.62" heatid="5003" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:26.91" heatid="23005" lane="2" />
                <ENTRY eventid="29" entrytime="00:02:43.55" heatid="29002" lane="4" />
                <ENTRY eventid="41" entrytime="00:05:11.62" heatid="41002" lane="4" />
                <ENTRY eventid="45" entrytime="00:00:00.00" heatid="45001" lane="3" />
                <ENTRY eventid="13" entrytime="00:01:10.87" heatid="13001" lane="7" />
                <ENTRY eventid="17" entrytime="00:01:22.77" heatid="17001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="62" eventid="1" swimtime="00:01:10.87" lane="6" heatid="1003" points="472" />
                <RESULT resultid="63" eventid="5" swimtime="00:01:22.77" lane="5" heatid="5003" points="465" />
                <RESULT resultid="808" eventid="13" swimtime="00:01:10.68" lane="7" heatid="13001" points="475" />
                <RESULT resultid="839" eventid="17" swimtime="00:01:19.85" lane="1" heatid="17001" points="518" />
                <RESULT resultid="64" eventid="23" swimtime="00:02:35.66" lane="2" heatid="23005" points="531">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="65" eventid="29" swimtime="00:02:47.25" lane="4" heatid="29002" points="556">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="66" eventid="41" swimtime="00:05:23.49" lane="4" heatid="41002" points="545">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.91" />
                    <SPLIT distance="200" swimtime="00:02:35.84" />
                    <SPLIT distance="300" swimtime="00:04:08.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="67" eventid="45" swimtime="00:04:53.27" lane="3" heatid="45001" points="517">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="200" swimtime="00:02:22.51" />
                    <SPLIT distance="300" swimtime="00:03:39.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="16" birthdate="2008-01-01" gender="M" lastname="Bodusch" firstname="Ben" license="377824" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:04.51" heatid="6002" lane="4" />
                <ENTRY eventid="22" entrytime="00:00:28.11" heatid="22003" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:25.98" heatid="28006" lane="3" />
                <ENTRY eventid="36" entrytime="00:00:57.58" heatid="36004" lane="4" />
                <ENTRY eventid="44" entrytime="00:00:31.07" heatid="44003" lane="3" />
                <ENTRY eventid="20" entrytime="00:01:10.44" heatid="20001" lane="5" />
                <ENTRY eventid="50" entrytime="00:01:04.62" heatid="50001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="68" eventid="6" swimtime="00:01:10.44" lane="4" heatid="6002" points="526" />
                <RESULT resultid="854" eventid="20" swimtime="00:01:08.34" lane="5" heatid="20001" points="576" />
                <RESULT resultid="69" eventid="22" swimtime="00:00:29.16" lane="3" heatid="22003" points="526" />
                <RESULT resultid="70" eventid="28" swimtime="00:00:26.30" lane="3" heatid="28006" points="607" />
                <RESULT resultid="71" eventid="36" swimtime="00:01:04.62" lane="4" heatid="36004" points="509" />
                <RESULT resultid="72" eventid="44" swimtime="00:00:31.24" lane="3" heatid="44003" points="573" />
                <RESULT resultid="911" eventid="50" swimtime="00:01:00.34" lane="3" heatid="50001" points="625" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="17" birthdate="2009-01-01" gender="F" lastname="Waizmann" firstname="Carlotta" license="391769" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:11.38" heatid="3003" lane="7" />
                <ENTRY eventid="11" entrytime="00:01:01.11" heatid="11005" lane="6" />
                <ENTRY eventid="21" entrytime="00:00:00.00" heatid="21001" lane="2" />
                <ENTRY eventid="35" entrytime="00:01:09.09" heatid="35005" lane="3" />
                <ENTRY eventid="39" entrytime="00:00:27.63" heatid="39004" lane="5" />
                <ENTRY eventid="32" entrytime="00:00:59.40" heatid="32001" lane="3" />
                <ENTRY eventid="48" entrytime="00:01:09.27" heatid="48001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="73" eventid="3" swimtime="00:02:08.90" lane="7" heatid="3003" points="660">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="74" eventid="11" swimtime="00:00:59.40" lane="6" heatid="11005" points="659" />
                <RESULT resultid="75" eventid="21" swimtime="00:00:31.76" lane="2" heatid="21001" points="604" />
                <RESULT resultid="866" eventid="32" swimtime="00:00:59.58" lane="3" heatid="32001" points="653" />
                <RESULT resultid="76" eventid="35" swimtime="00:01:09.27" lane="3" heatid="35005" points="560" />
                <RESULT resultid="77" eventid="39" swimtime="00:00:28.03" lane="5" heatid="39004" points="597" />
                <RESULT resultid="897" eventid="48" swimtime="00:01:08.53" lane="5" heatid="48001" points="579" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="18" birthdate="2012-01-01" gender="M" lastname="Severyuk" firstname="Daniel" license="440973" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:19.87" heatid="4002" lane="3" />
                <ENTRY eventid="8" entrytime="00:02:34.09" heatid="8002" lane="6" />
                <ENTRY eventid="24" entrytime="00:02:37.91" heatid="24002" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:28.82" heatid="28005" lane="2" />
                <ENTRY eventid="36" entrytime="00:01:12.36" heatid="36002" lane="7" />
                <ENTRY eventid="40" entrytime="00:00:29.35" heatid="40003" lane="7" />
                <ENTRY eventid="49" entrytime="00:01:08.15" heatid="49001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="78" eventid="4" swimtime="00:02:17.29" lane="3" heatid="4002" points="410">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="79" eventid="8" swimtime="00:02:32.35" lane="6" heatid="8002" points="396">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="80" eventid="24" swimtime="00:02:33.35" lane="3" heatid="24002" points="410">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="81" eventid="28" swimtime="00:00:29.44" lane="2" heatid="28005" points="432" />
                <RESULT resultid="82" eventid="36" swimtime="00:01:08.15" lane="7" heatid="36002" points="434" />
                <RESULT resultid="83" eventid="40" swimtime="00:00:28.74" lane="7" heatid="40003" points="385" />
                <RESULT resultid="905" eventid="49" swimtime="00:01:06.95" lane="2" heatid="49001" points="457" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="19" birthdate="2012-01-01" gender="F" lastname="Wießner" firstname="Emilia" license="434536" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:22.94" heatid="3002" lane="1" />
                <ENTRY eventid="11" entrytime="00:01:04.67" heatid="11003" lane="1" />
                <ENTRY eventid="23" entrytime="00:02:41.00" heatid="23003" lane="6" />
                <ENTRY eventid="27" entrytime="00:00:30.93" heatid="27004" lane="2" />
                <ENTRY eventid="39" entrytime="00:00:28.56" heatid="39003" lane="4" />
                <ENTRY eventid="45" entrytime="00:05:03.76" heatid="45003" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="84" eventid="3" swimtime="00:02:22.98" lane="1" heatid="3002" points="483">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="85" eventid="11" swimtime="00:01:04.56" lane="1" heatid="11003" points="513" />
                <RESULT resultid="86" eventid="23" swimtime="00:02:41.85" lane="6" heatid="23003" points="473">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="87" eventid="27" swimtime="00:00:31.76" lane="2" heatid="27004" points="455" />
                <RESULT resultid="88" eventid="39" swimtime="00:00:28.98" lane="4" heatid="39003" points="540" />
                <RESULT resultid="89" eventid="45" swimtime="00:05:09.38" lane="7" heatid="45003" points="440">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                    <SPLIT distance="200" swimtime="00:02:32.09" />
                    <SPLIT distance="300" swimtime="00:03:52.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="20" birthdate="2011-01-01" gender="F" lastname="Färber" firstname="Emma" license="408425" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:16.98" heatid="5002" lane="3" />
                <ENTRY eventid="11" entrytime="00:01:03.31" heatid="11003" lane="7" />
                <ENTRY eventid="21" entrytime="00:00:32.14" heatid="21003" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:31.08" heatid="27004" lane="7" />
                <ENTRY eventid="35" entrytime="00:01:10.11" heatid="35004" lane="6" />
                <ENTRY eventid="43" entrytime="00:00:40.10" heatid="43002" lane="7" />
                <ENTRY eventid="17" entrytime="00:01:19.10" heatid="17001" lane="6" />
                <ENTRY eventid="47" entrytime="00:01:11.46" heatid="47001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="90" eventid="5" swimtime="00:01:19.10" lane="3" heatid="5002" points="532" />
                <RESULT resultid="91" eventid="11" swimtime="00:01:04.59" lane="7" heatid="11003" points="513" />
                <RESULT resultid="836" eventid="17" swimtime="00:01:18.65" lane="6" heatid="17001" points="542" />
                <RESULT resultid="92" eventid="21" swimtime="00:00:33.55" lane="2" heatid="21003" points="513" />
                <RESULT resultid="93" eventid="27" status="DNS" swimtime="00:00:00.00" lane="7" heatid="27004" />
                <RESULT resultid="94" eventid="35" swimtime="00:01:11.46" lane="6" heatid="35004" points="510" />
                <RESULT resultid="95" eventid="43" swimtime="00:00:36.59" lane="7" heatid="43002" points="506" />
                <RESULT resultid="893" eventid="47" swimtime="00:01:09.53" lane="7" heatid="47001" points="554" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="21" birthdate="2013-01-01" gender="M" lastname="Brauer" firstname="Fabian" license="445392" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:09.54" heatid="2004" lane="1" />
                <ENTRY eventid="8" entrytime="00:02:38.92" heatid="8002" lane="7" />
                <ENTRY eventid="22" entrytime="00:00:34.60" heatid="22002" lane="4" />
                <ENTRY eventid="30" entrytime="00:03:06.53" heatid="30001" lane="3" />
                <ENTRY eventid="36" entrytime="00:01:16.82" heatid="36004" lane="8" />
                <ENTRY eventid="40" entrytime="00:00:29.09" heatid="40003" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="96" eventid="2" swimtime="00:01:08.80" lane="1" heatid="2004" points="371" />
                <RESULT resultid="97" eventid="8" swimtime="00:02:41.62" lane="7" heatid="8002" points="332">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="98" eventid="22" swimtime="00:00:33.57" lane="4" heatid="22002" points="345" />
                <RESULT resultid="99" eventid="30" swimtime="00:02:56.94" lane="3" heatid="30001" points="356">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="100" eventid="36" swimtime="00:01:12.49" lane="8" heatid="36004" points="360" />
                <RESULT resultid="101" eventid="40" swimtime="00:00:27.97" lane="2" heatid="40003" points="417" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="22" birthdate="2011-01-01" gender="M" lastname="Schoop" firstname="Finn" license="419064" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:06.57" heatid="2004" lane="7" />
                <ENTRY eventid="8" entrytime="00:02:25.53" heatid="8002" lane="5" />
                <ENTRY eventid="22" entrytime="00:00:30.04" heatid="22003" lane="2" />
                <ENTRY eventid="30" entrytime="00:02:45.27" heatid="30002" lane="1" />
                <ENTRY eventid="36" entrytime="00:01:05.71" heatid="36002" lane="3" />
                <ENTRY eventid="40" entrytime="00:00:27.51" heatid="40003" lane="4" />
                <ENTRY eventid="15" entrytime="00:01:05.18" heatid="15001" lane="6" />
                <ENTRY eventid="49" entrytime="00:01:05.34" heatid="49001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="102" eventid="2" swimtime="00:01:05.18" lane="7" heatid="2004" points="436" />
                <RESULT resultid="103" eventid="8" swimtime="00:02:23.67" lane="5" heatid="8002" points="472">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="821" eventid="15" swimtime="00:01:04.38" lane="6" heatid="15001" points="453" />
                <RESULT resultid="104" eventid="22" swimtime="00:00:29.90" lane="2" heatid="22003" points="488" />
                <RESULT resultid="105" eventid="30" swimtime="00:02:44.02" lane="1" heatid="30002" points="447">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="106" eventid="36" swimtime="00:01:05.34" lane="3" heatid="36002" points="492" />
                <RESULT resultid="107" eventid="40" swimtime="00:00:26.91" lane="4" heatid="40003" points="469" />
                <RESULT resultid="901" eventid="49" swimtime="00:01:04.42" lane="4" heatid="49001" points="513" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="23" birthdate="2005-01-01" gender="F" lastname="Vollmer" firstname="Hannah" license="341206" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:01.68" heatid="1004" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:28.07" heatid="27005" lane="4" />
                <ENTRY eventid="37" entrytime="00:02:15.84" heatid="37002" lane="4" />
                <ENTRY eventid="14" entrytime="00:01:05.26" heatid="14001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="108" eventid="1" swimtime="00:01:05.26" lane="4" heatid="1004" points="604" />
                <RESULT resultid="813" eventid="14" swimtime="00:01:04.58" lane="4" heatid="14001" points="623" />
                <RESULT resultid="109" eventid="27" swimtime="00:00:29.21" lane="4" heatid="27005" points="585" />
                <RESULT resultid="110" eventid="37" swimtime="00:02:29.37" lane="4" heatid="37002" points="542">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="24" birthdate="2011-01-01" gender="M" lastname="Frank" firstname="Hardy" license="423159" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:12.04" heatid="4003" lane="1" />
                <ENTRY eventid="12" entrytime="00:00:56.47" heatid="12005" lane="2" />
                <ENTRY eventid="24" entrytime="00:02:21.80" heatid="24004" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:29.31" heatid="28005" lane="1" />
                <ENTRY eventid="36" entrytime="00:01:10.34" heatid="36004" lane="7" />
                <ENTRY eventid="42" entrytime="00:05:25.29" heatid="42003" lane="2" />
                <ENTRY eventid="33" entrytime="00:00:58.05" heatid="33001" lane="6" />
                <ENTRY eventid="49" entrytime="00:01:08.90" heatid="49001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="111" eventid="4" swimtime="00:02:10.58" lane="1" heatid="4003" points="476">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="112" eventid="12" swimtime="00:00:58.05" lane="2" heatid="12005" points="510" />
                <RESULT resultid="113" eventid="24" swimtime="00:02:23.71" lane="1" heatid="24004" points="499">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="114" eventid="28" swimtime="00:00:28.09" lane="1" heatid="28005" points="498" />
                <RESULT resultid="874" eventid="33" swimtime="00:00:57.16" lane="6" heatid="33001" points="534" />
                <RESULT resultid="115" eventid="36" swimtime="00:01:08.90" lane="7" heatid="36004" points="420" />
                <RESULT resultid="116" eventid="42" swimtime="00:05:06.40" lane="2" heatid="42003" points="495">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="200" swimtime="00:02:31.03" />
                    <SPLIT distance="300" swimtime="00:03:58.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="907" eventid="49" swimtime="00:01:07.30" lane="1" heatid="49001" points="450" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="25" birthdate="2012-01-01" gender="F" lastname="Haupt" firstname="Helena Sophie" license="443234" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:24.67" heatid="5003" lane="2" />
                <ENTRY eventid="11" entrytime="00:01:03.05" heatid="11005" lane="7" />
                <ENTRY eventid="23" entrytime="00:02:38.10" heatid="23003" lane="5" />
                <ENTRY eventid="29" entrytime="00:03:11.86" heatid="29002" lane="8" />
                <ENTRY eventid="35" entrytime="00:01:13.36" heatid="35003" lane="7" />
                <ENTRY eventid="43" entrytime="00:00:38.88" heatid="43002" lane="5" />
                <ENTRY eventid="17" entrytime="00:01:23.51" heatid="17001" lane="8" />
                <ENTRY eventid="31" entrytime="00:01:03.75" heatid="31001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="117" eventid="5" swimtime="00:01:23.51" lane="2" heatid="5003" points="452" />
                <RESULT resultid="118" eventid="11" swimtime="00:01:03.75" lane="7" heatid="11005" points="533" />
                <RESULT resultid="840" eventid="17" swimtime="00:01:23.96" lane="8" heatid="17001" points="445" />
                <RESULT resultid="119" eventid="23" swimtime="00:02:36.21" lane="5" heatid="23003" points="526">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="120" eventid="29" swimtime="00:03:03.67" lane="8" heatid="29002" points="420">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="863" eventid="31" swimtime="00:01:06.16" lane="8" heatid="31001" points="477" />
                <RESULT resultid="121" eventid="35" swimtime="00:01:12.88" lane="7" heatid="35003" points="481" />
                <RESULT resultid="122" eventid="43" swimtime="00:00:37.78" lane="5" heatid="43002" points="459" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="26" birthdate="2010-01-01" gender="M" lastname="Harnisch" firstname="Henry" license="406011" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:05.71" heatid="4003" lane="3" />
                <ENTRY eventid="12" entrytime="00:00:57.08" heatid="12005" lane="7" />
                <ENTRY eventid="24" entrytime="00:02:20.32" heatid="24004" lane="7" />
                <ENTRY eventid="40" entrytime="00:00:26.74" heatid="40004" lane="6" />
                <ENTRY eventid="46" entrytime="00:04:21.89" heatid="46003" lane="6" />
                <ENTRY eventid="33" entrytime="00:00:57.73" heatid="33001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="123" eventid="4" swimtime="00:02:04.68" lane="3" heatid="4003" points="547">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="124" eventid="12" swimtime="00:00:57.73" lane="7" heatid="12005" points="519" />
                <RESULT resultid="125" eventid="24" swimtime="00:02:22.20" lane="7" heatid="24004" points="515">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="873" eventid="33" swimtime="00:00:57.82" lane="3" heatid="33001" points="516" />
                <RESULT resultid="126" eventid="40" swimtime="00:00:26.67" lane="6" heatid="40004" points="481" />
                <RESULT resultid="127" eventid="46" swimtime="00:04:24.73" lane="6" heatid="46003" points="574">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.52" />
                    <SPLIT distance="200" swimtime="00:02:09.74" />
                    <SPLIT distance="300" swimtime="00:03:17.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="27" birthdate="2007-01-01" gender="M" lastname="Reyher" firstname="Janek Thorben" license="361329" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:00.77" heatid="4004" lane="7" />
                <ENTRY eventid="12" entrytime="00:00:54.10" heatid="12003" lane="4" />
                <ENTRY eventid="22" entrytime="00:00:27.91" heatid="22003" lane="5" />
                <ENTRY eventid="30" entrytime="00:02:26.84" heatid="30002" lane="3" />
                <ENTRY eventid="40" entrytime="00:00:25.16" heatid="40005" lane="6" />
                <ENTRY eventid="44" entrytime="00:00:32.53" heatid="44003" lane="1" />
                <ENTRY eventid="34" entrytime="00:00:55.05" heatid="34001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="128" eventid="4" swimtime="00:01:59.03" lane="7" heatid="4004" points="629">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="129" eventid="12" swimtime="00:00:55.05" lane="4" heatid="12003" points="598" />
                <RESULT resultid="130" eventid="22" swimtime="00:00:28.30" lane="5" heatid="22003" points="576" />
                <RESULT resultid="131" eventid="30" swimtime="00:02:31.11" lane="3" heatid="30002" points="572">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="885" eventid="34" swimtime="00:00:57.40" lane="7" heatid="34001" points="528" />
                <RESULT resultid="132" eventid="40" swimtime="00:00:25.17" lane="6" heatid="40005" points="573" />
                <RESULT resultid="133" eventid="44" swimtime="00:00:32.76" lane="1" heatid="44003" points="497" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="28" birthdate="2007-01-01" gender="M" lastname="Herrmann" firstname="Jonas" license="366274" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:05.14" heatid="2005" lane="2" />
                <ENTRY eventid="8" entrytime="00:02:14.67" heatid="8003" lane="2" />
                <ENTRY eventid="24" entrytime="00:02:17.44" heatid="24004" lane="2" />
                <ENTRY eventid="36" entrytime="00:01:03.33" heatid="36003" lane="5" />
                <ENTRY eventid="40" entrytime="00:00:26.43" heatid="40004" lane="5" />
                <ENTRY eventid="16" entrytime="00:01:01.78" heatid="16001" lane="2" />
                <ENTRY eventid="50" entrytime="00:01:07.31" heatid="50001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="134" eventid="2" swimtime="00:01:01.78" lane="2" heatid="2005" points="512" />
                <RESULT resultid="135" eventid="8" swimtime="00:02:15.06" lane="2" heatid="8003" points="569">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="830" eventid="16" swimtime="00:01:01.39" lane="2" heatid="16001" points="522" />
                <RESULT resultid="136" eventid="24" swimtime="00:02:16.85" lane="2" heatid="24004" points="578">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="137" eventid="36" swimtime="00:01:07.31" lane="5" heatid="36003" points="450" />
                <RESULT resultid="138" eventid="40" swimtime="00:00:26.22" lane="5" heatid="40004" points="507" />
                <RESULT resultid="915" eventid="50" swimtime="00:01:03.56" lane="1" heatid="50001" points="535" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="29" birthdate="2013-01-01" gender="M" lastname="Richter" firstname="Justus" license="444299" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:24.75" heatid="6002" lane="6" />
                <ENTRY eventid="22" entrytime="00:00:36.88" heatid="22002" lane="2" />
                <ENTRY eventid="30" entrytime="00:02:57.17" heatid="30001" lane="5" />
                <ENTRY eventid="40" entrytime="00:00:31.51" heatid="40002" lane="1" />
                <ENTRY eventid="46" entrytime="00:05:06.48" heatid="46002" lane="7" />
                <ENTRY eventid="19" entrytime="00:01:25.10" heatid="19001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="139" eventid="6" swimtime="00:01:25.10" lane="6" heatid="6002" points="298" />
                <RESULT resultid="852" eventid="19" swimtime="00:01:24.49" lane="8" heatid="19001" points="305" />
                <RESULT resultid="140" eventid="22" swimtime="00:00:37.42" lane="2" heatid="22002" points="249" />
                <RESULT resultid="141" eventid="30" swimtime="00:02:57.18" lane="5" heatid="30001" points="355">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="142" eventid="40" swimtime="00:00:32.30" lane="1" heatid="40002" points="271" />
                <RESULT resultid="143" eventid="46" swimtime="00:05:12.42" lane="7" heatid="46002" points="349">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.46" />
                    <SPLIT distance="200" swimtime="00:02:34.69" />
                    <SPLIT distance="300" swimtime="00:03:55.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="30" birthdate="2009-01-01" gender="M" lastname="Baumeister" firstname="Lius Pepe" license="391171" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:00.92" heatid="2005" lane="3" />
                <ENTRY eventid="8" entrytime="00:02:12.36" heatid="8003" lane="6" />
                <ENTRY eventid="30" entrytime="00:02:27.63" heatid="30002" lane="6" />
                <ENTRY eventid="40" entrytime="00:00:26.13" heatid="40004" lane="4" />
                <ENTRY eventid="46" entrytime="00:04:09.30" heatid="46003" lane="5" />
                <ENTRY eventid="16" entrytime="00:01:01.33" heatid="16001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="144" eventid="2" swimtime="00:01:01.33" lane="3" heatid="2005" points="524" />
                <RESULT resultid="145" eventid="8" swimtime="00:02:12.69" lane="6" heatid="8003" points="600">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="829" eventid="16" swimtime="00:01:00.14" lane="6" heatid="16001" points="555" />
                <RESULT resultid="146" eventid="30" swimtime="00:02:26.33" lane="6" heatid="30002" points="630">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="147" eventid="40" swimtime="00:00:25.69" lane="4" heatid="40004" points="539" />
                <RESULT resultid="148" eventid="46" swimtime="00:04:10.89" lane="5" heatid="46003" points="674">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.10" />
                    <SPLIT distance="200" swimtime="00:02:02.57" />
                    <SPLIT distance="300" swimtime="00:03:06.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="31" birthdate="2004-01-01" gender="M" lastname="Schubert" firstname="Louis" license="358844" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:00:53.82" heatid="2005" lane="4" />
                <ENTRY eventid="12" entrytime="00:00:54.09" heatid="12004" lane="4" />
                <ENTRY eventid="38" entrytime="00:01:58.26" heatid="38002" lane="4" />
                <ENTRY eventid="40" entrytime="00:00:23.19" heatid="40005" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="149" eventid="2" status="WDR" swimtime="00:00:00.00" lane="4" heatid="2005" />
                <RESULT resultid="150" eventid="12" status="WDR" swimtime="00:00:00.00" lane="4" heatid="12004" />
                <RESULT resultid="151" eventid="38" status="WDR" swimtime="00:00:00.00" lane="4" heatid="38002" />
                <RESULT resultid="152" eventid="40" status="WDR" swimtime="00:00:00.00" lane="4" heatid="40005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="32" birthdate="2012-01-01" gender="F" lastname="Hacker" firstname="Mara" license="440971" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:15.83" heatid="1001" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:44.72" heatid="23002" lane="5" />
                <ENTRY eventid="27" entrytime="00:00:33.23" heatid="27003" lane="2" />
                <ENTRY eventid="37" entrytime="00:02:53.93" heatid="37002" lane="7" />
                <ENTRY eventid="43" entrytime="00:00:42.15" heatid="43001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="153" eventid="1" swimtime="00:01:13.51" lane="5" heatid="1001" points="422" />
                <RESULT resultid="154" eventid="23" swimtime="00:02:40.93" lane="5" heatid="23002" points="481">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="155" eventid="27" swimtime="00:00:32.50" lane="2" heatid="27003" points="424" />
                <RESULT resultid="156" eventid="37" swimtime="00:02:46.77" lane="7" heatid="37002" points="389">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="157" eventid="43" swimtime="00:00:39.18" lane="4" heatid="43001" points="412" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="33" birthdate="2009-01-01" gender="M" lastname="Jung" firstname="Marlon" license="391282" license_dbs="101860" license_dsv="391282" license_ipc="0" nation="GER">
              <HANDICAP free="S--" breast="SB--" medley="SM--" exception="12+" />
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:11.86" heatid="4003" lane="7" />
                <ENTRY eventid="10" entrytime="00:09:23.35" heatid="10000" lane="0" />
                <ENTRY eventid="24" entrytime="00:02:27.73" heatid="24003" lane="3" />
                <ENTRY eventid="30" entrytime="00:02:52.06" heatid="30001" lane="4" />
                <ENTRY eventid="42" entrytime="00:05:08.91" heatid="42000" lane="0" />
                <ENTRY eventid="46" entrytime="00:04:33.94" heatid="46000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="158" eventid="4" status="WDR" swimtime="00:00:00.00" lane="7" heatid="4003" />
                <RESULT resultid="159" eventid="10" status="WDR" swimtime="00:00:00.00" lane="0" heatid="10000" />
                <RESULT resultid="160" eventid="24" status="WDR" swimtime="00:00:00.00" lane="3" heatid="24003" />
                <RESULT resultid="161" eventid="30" status="WDR" swimtime="00:00:00.00" lane="4" heatid="30001" />
                <RESULT resultid="162" eventid="42" status="WDR" swimtime="00:00:00.00" lane="0" heatid="42000" />
                <RESULT resultid="163" eventid="46" status="WDR" swimtime="00:00:00.00" lane="0" heatid="46000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="34" birthdate="2008-01-01" gender="F" lastname="Rosenberg" firstname="Meike" license="373695" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:06.78" heatid="1002" lane="3" />
                <ENTRY eventid="7" entrytime="00:00:00.00" heatid="7001" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:00.00" heatid="27001" lane="3" />
                <ENTRY eventid="35" entrytime="00:00:00.00" heatid="35001" lane="7" />
                <ENTRY eventid="43" entrytime="00:00:36.07" heatid="43003" lane="2" />
                <ENTRY eventid="14" entrytime="00:01:06.61" heatid="14001" lane="2" />
                <ENTRY eventid="48" entrytime="00:01:09.79" heatid="48001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="164" eventid="1" swimtime="00:01:06.61" lane="3" heatid="1002" points="568" />
                <RESULT resultid="165" eventid="7" swimtime="00:02:31.00" lane="1" heatid="7001" points="542">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="817" eventid="14" swimtime="00:01:06.42" lane="2" heatid="14001" points="573" />
                <RESULT resultid="166" eventid="27" swimtime="00:00:29.32" lane="3" heatid="27001" points="578" />
                <RESULT resultid="167" eventid="35" swimtime="00:01:09.79" lane="7" heatid="35001" points="548" />
                <RESULT resultid="168" eventid="43" swimtime="00:00:36.83" lane="2" heatid="43003" points="496" />
                <RESULT resultid="899" eventid="48" swimtime="00:01:08.62" lane="6" heatid="48001" points="577" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="35" birthdate="2010-01-01" gender="F" lastname="Lißner" firstname="Mercedesz" license="426137" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:03.97" heatid="1003" lane="5" />
                <ENTRY eventid="5" entrytime="00:00:00.00" heatid="5003" lane="1" />
                <ENTRY eventid="11" entrytime="00:01:01.37" heatid="11004" lane="6" />
                <ENTRY eventid="27" entrytime="00:00:29.43" heatid="27005" lane="7" />
                <ENTRY eventid="39" entrytime="00:00:28.84" heatid="39003" lane="6" />
                <ENTRY eventid="45" entrytime="00:00:00.00" heatid="45001" lane="5" />
                <ENTRY eventid="13" entrytime="00:01:05.87" heatid="13001" lane="4" />
                <ENTRY eventid="17" entrytime="00:01:21.78" heatid="17001" lane="7" />
                <ENTRY eventid="31" entrytime="00:01:03.24" heatid="31001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="169" eventid="1" swimtime="00:01:05.87" lane="5" heatid="1003" points="587" />
                <RESULT resultid="170" eventid="5" swimtime="00:01:21.78" lane="1" heatid="5003" points="482" />
                <RESULT resultid="171" eventid="11" swimtime="00:01:03.24" lane="6" heatid="11004" points="546" />
                <RESULT resultid="803" eventid="13" swimtime="00:01:06.13" lane="4" heatid="13001" points="580" />
                <RESULT resultid="838" eventid="17" swimtime="00:01:20.97" lane="7" heatid="17001" points="496" />
                <RESULT resultid="172" eventid="27" swimtime="00:00:29.98" lane="7" heatid="27005" points="541" />
                <RESULT resultid="861" eventid="31" swimtime="00:01:03.28" lane="7" heatid="31001" points="545" />
                <RESULT resultid="173" eventid="39" swimtime="00:00:28.96" lane="6" heatid="39003" points="541" />
                <RESULT resultid="174" eventid="45" swimtime="00:04:47.69" lane="5" heatid="45001" points="547">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.74" />
                    <SPLIT distance="200" swimtime="00:02:18.43" />
                    <SPLIT distance="300" swimtime="00:03:33.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="36" birthdate="2012-01-01" gender="M" lastname="Birgel" firstname="Mick Günter" license="407310" nation="GER">
              <ENTRIES>
                <ENTRY eventid="8" entrytime="00:02:20.48" heatid="8002" lane="4" />
                <ENTRY eventid="12" entrytime="00:00:59.17" heatid="12003" lane="7" />
                <ENTRY eventid="24" entrytime="00:02:29.69" heatid="24003" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:29.52" heatid="28004" lane="4" />
                <ENTRY eventid="38" entrytime="00:02:37.56" heatid="38001" lane="4" />
                <ENTRY eventid="44" entrytime="00:00:38.64" heatid="44002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="175" eventid="8" swimtime="00:02:24.87" lane="4" heatid="8002" points="461">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="176" eventid="12" swimtime="00:01:00.20" lane="7" heatid="12003" points="457" />
                <RESULT resultid="177" eventid="24" swimtime="00:02:29.11" lane="1" heatid="24003" points="446">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="178" eventid="28" swimtime="00:00:29.29" lane="4" heatid="28004" points="439" />
                <RESULT resultid="179" eventid="38" swimtime="00:02:29.15" lane="4" heatid="38001" points="404">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="180" eventid="44" swimtime="00:00:37.44" lane="3" heatid="44002" points="332" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="37" birthdate="2008-01-01" gender="F" lastname="Clauß" firstname="Nele" license="366218" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:03.87" heatid="1004" lane="5" />
                <ENTRY eventid="7" entrytime="00:02:31.40" heatid="7002" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:33.39" heatid="23004" lane="3" />
                <ENTRY eventid="37" entrytime="00:02:21.63" heatid="37002" lane="3" />
                <ENTRY eventid="43" entrytime="00:00:38.95" heatid="43002" lane="3" />
                <ENTRY eventid="14" entrytime="00:01:06.24" heatid="14001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="181" eventid="1" swimtime="00:01:06.24" lane="5" heatid="1004" points="578" />
                <RESULT resultid="182" eventid="7" swimtime="00:02:35.08" lane="5" heatid="7002" points="500">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="815" eventid="14" swimtime="00:01:06.75" lane="3" heatid="14001" points="564" />
                <RESULT resultid="183" eventid="23" swimtime="00:02:35.55" lane="3" heatid="23004" points="533">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="184" eventid="37" swimtime="00:02:28.44" lane="3" heatid="37002" points="552">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="185" eventid="43" swimtime="00:00:39.75" lane="3" heatid="43002" points="394" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="38" birthdate="2010-01-01" gender="M" lastname="Turich" firstname="Niklas" license="417679" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:19.12" heatid="2002" lane="4" />
                <ENTRY eventid="8" entrytime="00:02:17.26" heatid="8003" lane="1" />
                <ENTRY eventid="24" entrytime="00:02:31.84" heatid="24003" lane="8" />
                <ENTRY eventid="40" entrytime="00:00:27.76" heatid="40003" lane="5" />
                <ENTRY eventid="46" entrytime="00:04:43.33" heatid="46003" lane="8" />
                <ENTRY eventid="15" entrytime="00:01:05.99" heatid="15001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="186" eventid="2" swimtime="00:01:05.99" lane="4" heatid="2002" points="420" />
                <RESULT resultid="187" eventid="8" swimtime="00:02:20.13" lane="1" heatid="8003" points="509">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="825" eventid="15" swimtime="00:01:04.59" lane="8" heatid="15001" points="448" />
                <RESULT resultid="188" eventid="24" swimtime="00:02:24.71" lane="8" heatid="24003" points="488">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="189" eventid="40" swimtime="00:00:26.80" lane="5" heatid="40003" points="474" />
                <RESULT resultid="190" eventid="46" swimtime="00:04:44.31" lane="8" heatid="46003" points="463">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="200" swimtime="00:02:20.18" />
                    <SPLIT distance="300" swimtime="00:03:32.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="39" birthdate="2011-01-01" gender="F" lastname="Schönberg" firstname="Ninett" license="418811" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:10.36" heatid="1003" lane="2" />
                <ENTRY eventid="11" entrytime="00:01:00.34" heatid="11003" lane="5" />
                <ENTRY eventid="23" entrytime="00:02:31.09" heatid="23005" lane="8" />
                <ENTRY eventid="35" entrytime="00:01:14.02" heatid="35003" lane="1" />
                <ENTRY eventid="39" entrytime="00:00:27.48" heatid="39005" lane="8" />
                <ENTRY eventid="13" entrytime="00:01:11.15" heatid="13001" lane="1" />
                <ENTRY eventid="31" entrytime="00:01:00.78" heatid="31001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="191" eventid="1" swimtime="00:01:11.15" lane="2" heatid="1003" points="466" />
                <RESULT resultid="192" eventid="11" swimtime="00:01:00.78" lane="5" heatid="11003" points="615" />
                <RESULT resultid="809" eventid="13" swimtime="00:01:11.15" lane="1" heatid="13001" points="466" />
                <RESULT resultid="193" eventid="23" swimtime="00:02:37.41" lane="8" heatid="23005" points="514">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="857" eventid="31" swimtime="00:01:01.28" lane="5" heatid="31001" points="600" />
                <RESULT resultid="194" eventid="35" status="WDR" swimtime="00:00:00.00" lane="1" heatid="35003" />
                <RESULT resultid="195" eventid="39" status="WDR" swimtime="00:00:00.00" lane="8" heatid="39005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="40" birthdate="2013-01-01" gender="F" lastname="Lißner" firstname="Phoebe" license="448337" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:12.85" heatid="1004" lane="1" />
                <ENTRY eventid="7" entrytime="00:02:34.23" heatid="7002" lane="2" />
                <ENTRY eventid="23" entrytime="00:02:36.49" heatid="23004" lane="1" />
                <ENTRY eventid="27" entrytime="00:00:32.44" heatid="27003" lane="6" />
                <ENTRY eventid="35" entrytime="00:01:11.42" heatid="35004" lane="2" />
                <ENTRY eventid="41" entrytime="00:05:43.99" heatid="41002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="196" eventid="1" swimtime="00:01:14.30" lane="1" heatid="1004" points="409" />
                <RESULT resultid="197" eventid="7" swimtime="00:02:40.58" lane="2" heatid="7002" points="450">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="198" eventid="23" swimtime="00:02:39.63" lane="1" heatid="23004" points="493">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="199" eventid="27" swimtime="00:00:31.84" lane="6" heatid="27003" points="451" />
                <RESULT resultid="200" eventid="35" swimtime="00:01:13.30" lane="2" heatid="35004" points="473" />
                <RESULT resultid="201" eventid="41" swimtime="00:05:40.54" lane="3" heatid="41002" points="467">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="200" swimtime="00:02:45.69" />
                    <SPLIT distance="300" swimtime="00:04:24.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="41" birthdate="2010-01-01" gender="F" lastname="Stodolka" firstname="Ronja" license="406010" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:10.48" heatid="1002" lane="2" />
                <ENTRY eventid="7" entrytime="00:00:00.00" heatid="7001" lane="7" />
                <ENTRY eventid="29" entrytime="00:02:47.78" heatid="29002" lane="3" />
                <ENTRY eventid="35" entrytime="00:01:16.32" heatid="35002" lane="4" />
                <ENTRY eventid="39" entrytime="00:00:00.00" heatid="39001" lane="6" />
                <ENTRY eventid="43" entrytime="00:00:36.12" heatid="43003" lane="7" />
                <ENTRY eventid="13" entrytime="00:01:11.47" heatid="13001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="202" eventid="1" swimtime="00:01:11.47" lane="2" heatid="1002" points="460" />
                <RESULT resultid="203" eventid="7" swimtime="00:02:34.68" lane="7" heatid="7001" points="504">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="810" eventid="13" swimtime="00:01:11.50" lane="8" heatid="13001" points="459" />
                <RESULT resultid="204" eventid="29" swimtime="00:02:47.63" lane="3" heatid="29002" points="552">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="205" eventid="35" swimtime="00:01:13.31" lane="4" heatid="35002" points="473" />
                <RESULT resultid="206" eventid="39" swimtime="00:00:30.09" lane="6" heatid="39001" points="483" />
                <RESULT resultid="207" eventid="43" swimtime="00:00:37.11" lane="7" heatid="43003" points="485" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="42" birthdate="2012-01-01" gender="F" lastname="Schindler" firstname="Rosa" license="440950" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:30.39" heatid="3001" lane="4" />
                <ENTRY eventid="9" entrytime="00:10:53.23" heatid="9002" lane="1" />
                <ENTRY eventid="21" entrytime="00:00:35.52" heatid="21002" lane="6" />
                <ENTRY eventid="27" entrytime="00:00:33.68" heatid="27003" lane="1" />
                <ENTRY eventid="39" entrytime="00:00:31.62" heatid="39002" lane="7" />
                <ENTRY eventid="45" entrytime="00:05:17.67" heatid="45002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="208" eventid="3" swimtime="00:02:28.97" lane="4" heatid="3001" points="427">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="209" eventid="9" swimtime="00:10:37.78" lane="1" heatid="9002" points="439">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="200" swimtime="00:02:34.86" />
                    <SPLIT distance="300" swimtime="00:03:54.80" />
                    <SPLIT distance="400" swimtime="00:05:15.68" />
                    <SPLIT distance="500" swimtime="00:06:37.25" />
                    <SPLIT distance="600" swimtime="00:07:58.67" />
                    <SPLIT distance="700" swimtime="00:09:20.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="210" eventid="21" swimtime="00:00:35.92" lane="6" heatid="21002" points="418" />
                <RESULT resultid="211" eventid="27" swimtime="00:00:33.00" lane="1" heatid="27003" points="405" />
                <RESULT resultid="212" eventid="39" swimtime="00:00:31.55" lane="7" heatid="39002" points="419" />
                <RESULT resultid="213" eventid="45" swimtime="00:05:11.86" lane="3" heatid="45002" points="429">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="200" swimtime="00:02:33.39" />
                    <SPLIT distance="300" swimtime="00:03:53.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="43" birthdate="2006-01-01" gender="F" lastname="Müller" firstname="Selina" license="349287" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:03.55" heatid="3003" lane="5" />
                <ENTRY eventid="11" entrytime="00:00:56.38" heatid="11005" lane="4" />
                <ENTRY eventid="25" entrytime="00:17:48.44" heatid="25001" lane="5" />
                <ENTRY eventid="39" entrytime="00:00:26.19" heatid="39005" lane="4" />
                <ENTRY eventid="32" entrytime="00:00:57.37" heatid="32001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="214" eventid="3" swimtime="00:02:05.90" lane="5" heatid="3003" points="708">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="215" eventid="11" swimtime="00:00:57.37" lane="4" heatid="11005" points="732" />
                <RESULT resultid="216" eventid="25" swimtime="00:17:32.69" lane="5" heatid="25001" points="668">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="200" swimtime="00:02:18.71" />
                    <SPLIT distance="300" swimtime="00:03:29.04" />
                    <SPLIT distance="400" swimtime="00:04:38.63" />
                    <SPLIT distance="500" swimtime="00:05:48.50" />
                    <SPLIT distance="600" swimtime="00:06:58.79" />
                    <SPLIT distance="700" swimtime="00:08:09.06" />
                    <SPLIT distance="800" swimtime="00:09:19.29" />
                    <SPLIT distance="900" swimtime="00:10:29.74" />
                    <SPLIT distance="1000" swimtime="00:11:41.13" />
                    <SPLIT distance="1100" swimtime="00:12:52.16" />
                    <SPLIT distance="1200" swimtime="00:14:03.16" />
                    <SPLIT distance="1300" swimtime="00:15:14.04" />
                    <SPLIT distance="1400" swimtime="00:16:24.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="864" eventid="32" swimtime="00:00:58.32" lane="4" heatid="32001" points="697" />
                <RESULT resultid="217" eventid="39" swimtime="00:00:26.69" lane="4" heatid="39005" points="692" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2008-01-01" gender="F" lastname="Luschnitz" firstname="Sophie" license="389677" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:11.94" heatid="3003" lane="1" />
                <ENTRY eventid="9" entrytime="00:09:35.14" heatid="9002" lane="3" />
                <ENTRY eventid="21" entrytime="00:00:00.00" heatid="21001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="218" eventid="3" swimtime="00:02:08.77" lane="1" heatid="3003" points="662">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="219" eventid="9" swimtime="00:09:35.85" lane="3" heatid="9002" points="596">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="200" swimtime="00:02:18.18" />
                    <SPLIT distance="300" swimtime="00:03:30.42" />
                    <SPLIT distance="400" swimtime="00:04:42.78" />
                    <SPLIT distance="500" swimtime="00:05:56.15" />
                    <SPLIT distance="600" swimtime="00:07:09.92" />
                    <SPLIT distance="700" swimtime="00:08:23.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="220" eventid="21" swimtime="00:00:31.60" lane="7" heatid="21001" points="614" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SSV 70 Halle-Neustadt" nation="GER" region="13" code="3603">
          <ATHLETES>
            <ATHLETE athleteid="66" birthdate="2014-01-01" gender="F" lastname="Schulz" firstname="Emma Leni" license="450929" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:43.84" heatid="3001" lane="2" />
                <ENTRY eventid="11" entrytime="00:01:14.77" heatid="11001" lane="4" />
                <ENTRY eventid="21" entrytime="00:00:37.22" heatid="21002" lane="1" />
                <ENTRY eventid="23" entrytime="00:02:54.83" heatid="23001" lane="3" />
                <ENTRY eventid="39" entrytime="00:00:33.36" heatid="39001" lane="4" />
                <ENTRY eventid="45" entrytime="00:05:42.72" heatid="45002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="315" eventid="3" swimtime="00:02:36.08" lane="2" heatid="3001" points="371">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="316" eventid="11" swimtime="00:01:10.91" lane="4" heatid="11001" points="387" />
                <RESULT resultid="317" eventid="21" swimtime="00:00:36.81" lane="1" heatid="21002" points="388" />
                <RESULT resultid="318" eventid="23" swimtime="00:02:59.25" lane="3" heatid="23001" points="348">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="319" eventid="39" swimtime="00:00:32.44" lane="4" heatid="39001" points="385" />
                <RESULT resultid="320" eventid="45" swimtime="00:05:27.62" lane="1" heatid="45002" points="370">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="200" swimtime="00:02:39.92" />
                    <SPLIT distance="300" swimtime="00:04:04.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="67" birthdate="2013-01-01" gender="M" lastname="Zorn" firstname="Jannik" license="450934" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:55.89" heatid="4001" lane="5" />
                <ENTRY eventid="12" entrytime="00:01:19.29" heatid="12001" lane="1" />
                <ENTRY eventid="24" entrytime="00:02:56.53" heatid="24001" lane="6" />
                <ENTRY eventid="28" entrytime="00:00:38.74" heatid="28002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="321" eventid="4" swimtime="00:02:39.27" lane="5" heatid="4001" points="262">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="322" eventid="12" swimtime="00:01:12.95" lane="1" heatid="12001" points="257" />
                <RESULT resultid="323" eventid="24" swimtime="00:02:52.43" lane="6" heatid="24001" points="288">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="324" eventid="28" swimtime="00:00:36.97" lane="1" heatid="28002" points="218" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="68" birthdate="2013-01-01" gender="F" lastname="Petzold" firstname="Luzie" license="450925" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:46.53" heatid="3001" lane="7" />
                <ENTRY eventid="11" entrytime="00:01:14.19" heatid="11002" lane="2" />
                <ENTRY eventid="23" entrytime="00:03:08.82" heatid="23001" lane="8" />
                <ENTRY eventid="27" entrytime="00:00:38.64" heatid="27001" lane="4" />
                <ENTRY eventid="35" entrytime="00:01:27.92" heatid="35001" lane="4" />
                <ENTRY eventid="45" entrytime="00:05:57.05" heatid="45001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="325" eventid="3" swimtime="00:02:47.71" lane="7" heatid="3001" points="299">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="326" eventid="11" swimtime="00:01:14.81" lane="2" heatid="11002" points="330" />
                <RESULT resultid="327" eventid="23" status="WDR" swimtime="00:00:00.00" lane="8" heatid="23001" />
                <RESULT resultid="328" eventid="27" status="WDR" swimtime="00:00:00.00" lane="4" heatid="27001" />
                <RESULT resultid="329" eventid="35" status="WDR" swimtime="00:00:00.00" lane="4" heatid="35001" />
                <RESULT resultid="330" eventid="45" status="WDR" swimtime="00:00:00.00" lane="4" heatid="45001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SSV Leutzsch" nation="GER" region="12" code="3378">
          <ATHLETES>
            <ATHLETE athleteid="158" birthdate="2004-01-01" gender="M" lastname="Vielland" firstname="Edwin" license="340594" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:03.83" heatid="2005" lane="6" />
                <ENTRY eventid="10" entrytime="00:09:20.00" heatid="10002" lane="6" />
                <ENTRY eventid="28" entrytime="00:00:29.65" heatid="28004" lane="5" />
                <ENTRY eventid="16" entrytime="00:01:04.07" heatid="16001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="737" eventid="2" swimtime="00:01:04.07" lane="6" heatid="2005" points="459" />
                <RESULT resultid="738" eventid="10" swimtime="00:09:29.98" lane="6" heatid="10002" points="499">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.25" />
                    <SPLIT distance="200" swimtime="00:02:14.01" />
                    <SPLIT distance="300" swimtime="00:03:25.46" />
                    <SPLIT distance="400" swimtime="00:04:38.18" />
                    <SPLIT distance="500" swimtime="00:05:51.48" />
                    <SPLIT distance="600" swimtime="00:07:05.02" />
                    <SPLIT distance="700" swimtime="00:08:18.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="832" eventid="16" swimtime="00:01:05.93" lane="1" heatid="16001" points="421" />
                <RESULT resultid="739" eventid="28" swimtime="00:00:29.32" lane="5" heatid="28004" points="438" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="159" birthdate="2006-01-01" gender="M" lastname="Plewa" firstname="Florian" license="345830" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:00.50" heatid="2003" lane="5" />
                <ENTRY eventid="12" entrytime="00:00:54.69" heatid="12004" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:26.39" heatid="28006" lane="6" />
                <ENTRY eventid="40" entrytime="00:00:25.44" heatid="40005" lane="2" />
                <ENTRY eventid="44" entrytime="00:00:32.50" heatid="44003" lane="7" />
                <ENTRY eventid="16" entrytime="00:00:59.25" heatid="16001" lane="5" />
                <ENTRY eventid="34" entrytime="00:00:54.83" heatid="34001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="740" eventid="2" swimtime="00:00:59.25" lane="5" heatid="2003" points="581" />
                <RESULT resultid="741" eventid="12" swimtime="00:00:54.83" lane="3" heatid="12004" points="606" />
                <RESULT resultid="827" eventid="16" swimtime="00:00:59.03" lane="5" heatid="16001" points="587" />
                <RESULT resultid="742" eventid="28" swimtime="00:00:25.93" lane="6" heatid="28006" points="633" />
                <RESULT resultid="883" eventid="34" swimtime="00:00:54.97" lane="6" heatid="34001" points="601" />
                <RESULT resultid="743" eventid="40" swimtime="00:00:24.63" lane="2" heatid="40005" points="611" />
                <RESULT resultid="744" eventid="44" swimtime="00:00:32.04" lane="7" heatid="44003" points="531" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2010-01-01" gender="M" lastname="Plewa" firstname="Richard" license="433622" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:04.10" heatid="2004" lane="6" />
                <ENTRY eventid="12" entrytime="00:01:00.65" heatid="12002" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:29.44" heatid="28005" lane="8" />
                <ENTRY eventid="40" entrytime="00:00:27.77" heatid="40003" lane="3" />
                <ENTRY eventid="44" entrytime="00:00:38.10" heatid="44002" lane="5" />
                <ENTRY eventid="15" entrytime="00:01:03.64" heatid="15001" lane="5" />
                <ENTRY eventid="33" entrytime="00:00:59.71" heatid="33001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="745" eventid="2" swimtime="00:01:03.64" lane="6" heatid="2004" points="469" />
                <RESULT resultid="746" eventid="12" swimtime="00:00:59.71" lane="4" heatid="12002" points="469" />
                <RESULT resultid="819" eventid="15" swimtime="00:01:02.56" lane="5" heatid="15001" points="493" />
                <RESULT resultid="747" eventid="28" swimtime="00:00:28.34" lane="8" heatid="28005" points="485" />
                <RESULT resultid="877" eventid="33" swimtime="00:00:59.97" lane="1" heatid="33001" points="463" />
                <RESULT resultid="748" eventid="40" swimtime="00:00:27.21" lane="3" heatid="40003" points="453" />
                <RESULT resultid="749" eventid="44" swimtime="00:00:36.36" lane="5" heatid="44002" points="363" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2013-01-01" gender="M" lastname="Plewa" firstname="Valentin" license="441003" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:20.34" heatid="2002" lane="5" />
                <ENTRY eventid="12" entrytime="00:01:10.26" heatid="12001" lane="5" />
                <ENTRY eventid="22" entrytime="00:00:37.75" heatid="22002" lane="7" />
                <ENTRY eventid="28" entrytime="00:00:32.73" heatid="28003" lane="6" />
                <ENTRY eventid="40" entrytime="00:00:30.60" heatid="40002" lane="6" />
                <ENTRY eventid="44" entrytime="00:00:42.71" heatid="44001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="750" eventid="2" swimtime="00:01:14.61" lane="5" heatid="2002" points="291" />
                <RESULT resultid="751" eventid="12" swimtime="00:01:08.90" lane="5" heatid="12001" points="305" />
                <RESULT resultid="752" eventid="22" swimtime="00:00:37.17" lane="7" heatid="22002" points="254" />
                <RESULT resultid="753" eventid="28" swimtime="00:00:32.82" lane="6" heatid="28003" points="312" />
                <RESULT resultid="754" eventid="40" swimtime="00:00:29.84" lane="6" heatid="40002" points="344" />
                <RESULT resultid="755" eventid="44" swimtime="00:00:39.70" lane="4" heatid="44001" points="279" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="ST Erzgebirge" nation="GER" region="12" code="5134">
          <ATHLETES>
            <ATHLETE athleteid="90" birthdate="2011-01-01" gender="F" lastname="Schreiter" firstname="Melissa" license="447078" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:23.49" heatid="5002" lane="6" />
                <ENTRY eventid="23" entrytime="00:02:43.50" heatid="23003" lane="7" />
                <ENTRY eventid="29" entrytime="00:02:58.50" heatid="29002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="434" eventid="5" swimtime="00:01:24.05" lane="6" heatid="5002" points="444" />
                <RESULT resultid="435" eventid="23" swimtime="00:02:42.17" lane="7" heatid="23003" points="470">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="436" eventid="29" swimtime="00:02:53.04" lane="2" heatid="29002" points="502">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="STV Limbach-Oberfrohna e.V." nation="GER" region="12" code="5406">
          <ATHLETES>
            <ATHLETE athleteid="157" birthdate="2007-01-01" gender="M" lastname="Straßburger" firstname="Christoph" license="349627" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:01:56.48" heatid="4004" lane="3" />
                <ENTRY eventid="12" entrytime="00:00:54.28" heatid="12004" lane="5" />
                <ENTRY eventid="38" entrytime="00:02:06.02" heatid="38002" lane="3" />
                <ENTRY eventid="34" entrytime="00:00:54.46" heatid="34001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="734" eventid="4" swimtime="00:01:57.90" lane="3" heatid="4004" points="647">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="735" eventid="12" swimtime="00:00:54.46" lane="5" heatid="12004" points="618" />
                <RESULT resultid="882" eventid="34" swimtime="00:00:54.52" lane="3" heatid="34001" points="616" />
                <RESULT resultid="736" eventid="38" swimtime="00:02:10.21" lane="3" heatid="38002" points="608">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV 1919 Grimma" nation="GER" region="12" code="5149">
          <ATHLETES>
            <ATHLETE athleteid="1" birthdate="2013-01-01" gender="M" lastname="Munari" firstname="Alessandro" license="445022" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:11:17.27" heatid="10001" lane="1" />
                <ENTRY eventid="24" entrytime="00:02:55.15" heatid="24001" lane="5" />
                <ENTRY eventid="40" entrytime="00:00:32.42" heatid="40001" lane="3" />
                <ENTRY eventid="46" entrytime="00:05:18.50" heatid="46002" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="1" eventid="10" swimtime="00:11:07.82" lane="1" heatid="10001" points="310">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.03" />
                    <SPLIT distance="200" swimtime="00:02:40.71" />
                    <SPLIT distance="300" swimtime="00:04:05.24" />
                    <SPLIT distance="400" swimtime="00:05:30.58" />
                    <SPLIT distance="500" swimtime="00:06:55.45" />
                    <SPLIT distance="600" swimtime="00:08:20.19" />
                    <SPLIT distance="700" swimtime="00:09:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2" eventid="24" swimtime="00:02:58.21" lane="5" heatid="24001" points="261">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3" eventid="40" swimtime="00:00:32.90" lane="3" heatid="40001" points="256" />
                <RESULT resultid="4" eventid="46" swimtime="00:05:19.58" lane="8" heatid="46002" points="326">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.85" />
                    <SPLIT distance="200" swimtime="00:02:36.70" />
                    <SPLIT distance="300" swimtime="00:03:58.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="2" birthdate="2005-01-01" gender="M" lastname="von Thun" firstname="Karl" license="329642" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:08:28.73" heatid="10002" lane="4" />
                <ENTRY eventid="28" entrytime="00:00:25.64" heatid="28006" lane="4" />
                <ENTRY eventid="38" entrytime="00:02:01.56" heatid="38002" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="5" eventid="10" swimtime="00:08:32.67" lane="4" heatid="10002" points="685">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.09" />
                    <SPLIT distance="200" swimtime="00:02:05.03" />
                    <SPLIT distance="300" swimtime="00:03:09.47" />
                    <SPLIT distance="400" swimtime="00:04:14.12" />
                    <SPLIT distance="500" swimtime="00:05:18.91" />
                    <SPLIT distance="600" swimtime="00:06:24.13" />
                    <SPLIT distance="700" swimtime="00:07:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6" eventid="28" swimtime="00:00:26.40" lane="4" heatid="28006" points="600" />
                <RESULT resultid="7" eventid="38" swimtime="00:02:06.35" lane="5" heatid="38002" points="665">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Halle / Saale" nation="GER" region="13" code="3593">
          <ATHLETES>
            <ATHLETE athleteid="91" birthdate="2011-01-01" gender="F" lastname="Hennig" firstname="Alice" license="420404" nation="GER">
              <ENTRIES>
                <ENTRY eventid="7" entrytime="00:02:26.47" heatid="7002" lane="4" />
                <ENTRY eventid="11" entrytime="00:00:59.89" heatid="11004" lane="5" />
                <ENTRY eventid="21" entrytime="00:00:31.90" heatid="21003" lane="3" />
                <ENTRY eventid="35" entrytime="00:01:07.59" heatid="35005" lane="5" />
                <ENTRY eventid="31" entrytime="00:01:00.87" heatid="31001" lane="3" />
                <ENTRY eventid="47" entrytime="00:01:10.16" heatid="47001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="437" eventid="7" swimtime="00:02:30.31" lane="4" heatid="7002" points="549">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="438" eventid="11" swimtime="00:01:00.87" lane="5" heatid="11004" points="613" />
                <RESULT resultid="439" eventid="21" swimtime="00:00:32.59" lane="3" heatid="21003" points="559" />
                <RESULT resultid="858" eventid="31" swimtime="00:01:01.12" lane="3" heatid="31001" points="605" />
                <RESULT resultid="440" eventid="35" swimtime="00:01:10.16" lane="5" heatid="35005" points="539" />
                <RESULT resultid="890" eventid="47" swimtime="00:01:10.57" lane="3" heatid="47001" points="530" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="92" birthdate="2010-01-01" gender="M" lastname="Riß" firstname="Bjarne" license="407283" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:05.73" heatid="2003" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:30.36" heatid="28004" lane="3" />
                <ENTRY eventid="38" entrytime="00:02:34.18" heatid="38002" lane="8" />
                <ENTRY eventid="15" entrytime="00:01:05.31" heatid="15001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="441" eventid="2" swimtime="00:01:05.31" lane="2" heatid="2003" points="434" />
                <RESULT resultid="823" eventid="15" swimtime="00:01:05.52" lane="7" heatid="15001" points="429" />
                <RESULT resultid="442" eventid="28" swimtime="00:00:29.38" lane="3" heatid="28004" points="435" />
                <RESULT resultid="443" eventid="38" swimtime="00:02:29.72" lane="8" heatid="38002" points="400">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="93" birthdate="2011-01-01" gender="M" lastname="Waletzki" firstname="Bruno" license="427152" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:08.29" heatid="4003" lane="6" />
                <ENTRY eventid="12" entrytime="00:00:55.85" heatid="12005" lane="6" />
                <ENTRY eventid="36" entrytime="00:01:09.19" heatid="36002" lane="2" />
                <ENTRY eventid="33" entrytime="00:00:55.97" heatid="33001" lane="4" />
                <ENTRY eventid="49" entrytime="00:01:06.91" heatid="49001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="444" eventid="4" swimtime="00:02:04.39" lane="6" heatid="4003" points="551">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="445" eventid="12" swimtime="00:00:55.97" lane="6" heatid="12005" points="569" />
                <RESULT resultid="871" eventid="33" swimtime="00:00:56.00" lane="4" heatid="33001" points="568" />
                <RESULT resultid="446" eventid="36" swimtime="00:01:06.91" lane="2" heatid="36002" points="458" />
                <RESULT resultid="903" eventid="49" swimtime="00:01:06.77" lane="3" heatid="49001" points="461" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="94" birthdate="2008-01-01" gender="F" lastname="Klemm" firstname="Charlotte Maria" license="402158">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:11.34" heatid="3003" lane="2" />
                <ENTRY eventid="23" entrytime="00:02:20.96" heatid="23005" lane="5" />
                <ENTRY eventid="39" entrytime="00:00:26.98" heatid="39005" lane="5" />
                <ENTRY eventid="43" entrytime="00:00:33.01" heatid="43003" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="447" eventid="3" swimtime="00:02:08.13" lane="2" heatid="3003" points="672">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="448" eventid="23" swimtime="00:02:20.92" lane="5" heatid="23005" points="716">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="449" eventid="39" swimtime="00:00:27.28" lane="5" heatid="39005" points="648" />
                <RESULT resultid="450" eventid="43" swimtime="00:00:34.26" lane="4" heatid="43003" points="616" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="95" birthdate="2008-01-01" gender="M" lastname="Stark" firstname="Clemens" license="379642" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:01.16" heatid="4004" lane="8" />
                <ENTRY eventid="12" entrytime="00:00:54.54" heatid="12005" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:28.87" heatid="28005" lane="7" />
                <ENTRY eventid="40" entrytime="00:00:24.34" heatid="40005" lane="5" />
                <ENTRY eventid="34" entrytime="00:00:55.48" heatid="34000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="451" eventid="4" swimtime="00:02:07.37" lane="8" heatid="4004" points="513">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="452" eventid="12" swimtime="00:00:55.48" lane="3" heatid="12005" points="584" />
                <RESULT resultid="453" eventid="28" status="DNS" swimtime="00:00:00.00" lane="7" heatid="28005" />
                <RESULT resultid="879" eventid="34" status="WDR" swimtime="00:00:00.00" lane="0" heatid="34000" />
                <RESULT resultid="454" eventid="40" swimtime="00:00:24.55" lane="5" heatid="40005" points="617" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="96" birthdate="2010-01-01" gender="M" lastname="Prade" firstname="Dominik" license="414210" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:05.26" heatid="2004" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:28.70" heatid="28005" lane="6" />
                <ENTRY eventid="38" entrytime="00:02:20.58" heatid="38002" lane="7" />
                <ENTRY eventid="44" entrytime="00:00:38.91" heatid="44002" lane="6" />
                <ENTRY eventid="15" entrytime="00:01:03.72" heatid="15001" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="455" eventid="2" swimtime="00:01:03.72" lane="2" heatid="2004" points="467" />
                <RESULT resultid="820" eventid="15" swimtime="00:01:03.42" lane="3" heatid="15001" points="474" />
                <RESULT resultid="456" eventid="28" swimtime="00:00:28.27" lane="6" heatid="28005" points="488" />
                <RESULT resultid="457" eventid="38" swimtime="00:02:25.28" lane="7" heatid="38002" points="438">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="458" eventid="44" swimtime="00:00:37.17" lane="6" heatid="44002" points="340" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="97" birthdate="2009-01-01" gender="M" lastname="Böhme" firstname="Erik Sebastian" license="409018" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:08.67" heatid="4000" lane="0" />
                <ENTRY eventid="24" entrytime="00:02:24.76" heatid="24000" lane="0" />
                <ENTRY eventid="40" entrytime="00:00:29.21" heatid="40000" lane="0" />
                <ENTRY eventid="44" entrytime="00:00:40.63" heatid="44000" lane="0" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="459" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="460" eventid="24" status="WDR" swimtime="00:00:00.00" lane="0" heatid="24000" />
                <RESULT resultid="461" eventid="40" status="WDR" swimtime="00:00:00.00" lane="0" heatid="40000" />
                <RESULT resultid="462" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="98" birthdate="2010-01-01" gender="F" lastname="Hilbich" firstname="Fiona Sophie" license="419502" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:16.64" heatid="5001" lane="5" />
                <ENTRY eventid="27" entrytime="00:00:31.13" heatid="27004" lane="1" />
                <ENTRY eventid="39" entrytime="00:00:30.83" heatid="39002" lane="2" />
                <ENTRY eventid="43" entrytime="00:00:36.70" heatid="43003" lane="1" />
                <ENTRY eventid="17" entrytime="00:01:17.84" heatid="17001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="463" eventid="5" swimtime="00:01:17.84" lane="5" heatid="5001" points="559" />
                <RESULT resultid="833" eventid="17" swimtime="00:01:17.79" lane="4" heatid="17001" points="560" />
                <RESULT resultid="464" eventid="27" swimtime="00:00:31.46" lane="1" heatid="27004" points="468" />
                <RESULT resultid="465" eventid="39" swimtime="00:00:29.20" lane="2" heatid="39002" points="528" />
                <RESULT resultid="466" eventid="43" swimtime="00:00:38.26" lane="1" heatid="43003" points="442" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="99" birthdate="2007-01-01" gender="M" lastname="Leineweber" firstname="Florian Paul" license="337373" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:05.00" heatid="4003" lane="5" />
                <ENTRY eventid="12" entrytime="00:01:00.00" heatid="12003" lane="1" />
                <ENTRY eventid="40" entrytime="00:00:25.00" heatid="40005" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="467" eventid="4" swimtime="00:02:05.07" lane="5" heatid="4003" points="542">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="468" eventid="12" swimtime="00:00:58.00" lane="1" heatid="12003" points="512" />
                <RESULT resultid="469" eventid="40" swimtime="00:00:26.18" lane="3" heatid="40005" points="509" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100" birthdate="2012-01-01" gender="M" lastname="Tanke" firstname="Fynn Valentin" license="448146" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:09:55.00" heatid="10001" lane="4" />
                <ENTRY eventid="24" entrytime="00:02:29.13" heatid="24003" lane="7" />
                <ENTRY eventid="42" entrytime="00:05:38.85" heatid="42003" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="470" eventid="10" swimtime="00:09:38.81" lane="4" heatid="10001" points="476">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.61" />
                    <SPLIT distance="200" swimtime="00:02:18.76" />
                    <SPLIT distance="300" swimtime="00:03:32.39" />
                    <SPLIT distance="400" swimtime="00:04:46.95" />
                    <SPLIT distance="500" swimtime="00:06:01.14" />
                    <SPLIT distance="600" swimtime="00:07:15.25" />
                    <SPLIT distance="700" swimtime="00:08:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="471" eventid="24" swimtime="00:02:29.10" lane="7" heatid="24003" points="446">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="472" eventid="42" swimtime="00:05:20.38" lane="8" heatid="42003" points="433">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.21" />
                    <SPLIT distance="200" swimtime="00:02:36.89" />
                    <SPLIT distance="300" swimtime="00:04:09.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101" birthdate="2010-01-01" gender="M" lastname="Schenk" firstname="Georg Maximilian" license="429218" nation="GER">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:11.26" heatid="6003" lane="5" />
                <ENTRY eventid="30" entrytime="00:02:34.88" heatid="30002" lane="2" />
                <ENTRY eventid="42" entrytime="00:05:05.42" heatid="42003" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:14.20" heatid="19001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="473" eventid="6" swimtime="00:01:14.20" lane="5" heatid="6003" points="450" />
                <RESULT resultid="846" eventid="19" swimtime="00:01:12.83" lane="5" heatid="19001" points="476" />
                <RESULT resultid="474" eventid="30" swimtime="00:02:38.77" lane="2" heatid="30002" points="493">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="475" eventid="42" swimtime="00:05:12.13" lane="4" heatid="42003" points="468">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.39" />
                    <SPLIT distance="200" swimtime="00:02:31.39" />
                    <SPLIT distance="300" swimtime="00:04:00.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102" birthdate="2012-01-01" gender="F" lastname="Erhard" firstname="Ida" license="426571" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:13.69" heatid="1003" lane="1" />
                <ENTRY eventid="9" entrytime="00:11:18.94" heatid="9002" lane="8" />
                <ENTRY eventid="21" entrytime="00:00:34.91" heatid="21002" lane="3" />
                <ENTRY eventid="23" entrytime="00:02:44.14" heatid="23003" lane="1" />
                <ENTRY eventid="41" entrytime="00:06:19.04" heatid="41002" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="476" eventid="1" swimtime="00:01:12.36" lane="1" heatid="1003" points="443" />
                <RESULT resultid="477" eventid="9" swimtime="00:10:25.25" lane="8" heatid="9002" points="466">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.48" />
                    <SPLIT distance="200" swimtime="00:02:33.57" />
                    <SPLIT distance="300" swimtime="00:03:52.89" />
                    <SPLIT distance="400" swimtime="00:05:12.63" />
                    <SPLIT distance="500" swimtime="00:06:32.22" />
                    <SPLIT distance="600" swimtime="00:07:51.13" />
                    <SPLIT distance="700" swimtime="00:09:10.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="478" eventid="21" swimtime="00:00:35.94" lane="3" heatid="21002" points="417" />
                <RESULT resultid="479" eventid="23" swimtime="00:02:43.24" lane="1" heatid="23003" points="461">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="480" eventid="41" swimtime="00:05:42.57" lane="1" heatid="41002" points="459">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.69" />
                    <SPLIT distance="200" swimtime="00:02:41.40" />
                    <SPLIT distance="300" swimtime="00:04:28.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="103" birthdate="2011-01-01" gender="M" lastname="Stark" firstname="Jakob" license="413607">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:15.59" heatid="4003" lane="8" />
                <ENTRY eventid="12" entrytime="00:01:01.68" heatid="12002" lane="5" />
                <ENTRY eventid="22" entrytime="00:00:30.00" heatid="22003" lane="6" />
                <ENTRY eventid="42" entrytime="00:05:26.99" heatid="42003" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="481" eventid="4" swimtime="00:02:14.69" lane="8" heatid="4003" points="434">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="482" eventid="12" swimtime="00:00:59.95" lane="5" heatid="12002" points="463" />
                <RESULT resultid="483" eventid="22" swimtime="00:00:35.40" lane="6" heatid="22003" points="294" />
                <RESULT resultid="484" eventid="42" swimtime="00:05:21.67" lane="7" heatid="42003" points="428">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="200" swimtime="00:02:41.61" />
                    <SPLIT distance="300" swimtime="00:04:10.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="104" birthdate="2014-01-01" gender="M" lastname="Jäger" firstname="Jan" license="450452" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:53.47" heatid="4001" lane="4" />
                <ENTRY eventid="8" entrytime="00:03:14.41" heatid="8001" lane="3" />
                <ENTRY eventid="24" entrytime="00:03:13.33" heatid="24001" lane="1" />
                <ENTRY eventid="28" entrytime="00:00:38.60" heatid="28002" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="485" eventid="4" swimtime="00:02:40.62" lane="4" heatid="4001" points="256">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="486" eventid="8" swimtime="00:03:12.56" lane="3" heatid="8001" points="196">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="487" eventid="24" swimtime="00:03:11.69" lane="1" heatid="24001" points="210">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="488" eventid="28" swimtime="00:00:37.57" lane="7" heatid="28002" points="208" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105" birthdate="2005-01-01" gender="M" lastname="Bohnert" firstname="Jules" license="339244" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:00:55.86" heatid="2004" lane="4" />
                <ENTRY eventid="12" entrytime="00:00:54.53" heatid="12003" lane="5" />
                <ENTRY eventid="28" entrytime="00:00:25.83" heatid="28006" lane="5" />
                <ENTRY eventid="16" entrytime="00:00:56.31" heatid="16001" lane="4" />
                <ENTRY eventid="34" entrytime="00:00:53.06" heatid="34001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="489" eventid="2" swimtime="00:00:56.31" lane="4" heatid="2004" points="677" />
                <RESULT resultid="490" eventid="12" swimtime="00:00:53.06" lane="5" heatid="12003" points="668" />
                <RESULT resultid="826" eventid="16" swimtime="00:00:56.69" lane="4" heatid="16001" points="663" />
                <RESULT resultid="491" eventid="28" swimtime="00:00:27.74" lane="5" heatid="28006" points="517" />
                <RESULT resultid="880" eventid="34" swimtime="00:00:53.61" lane="4" heatid="34001" points="648" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106" birthdate="2006-01-01" gender="F" lastname="Heinze" firstname="Juliane" license="356548">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:04.77" heatid="1004" lane="3" />
                <ENTRY eventid="11" entrytime="00:00:59.41" heatid="11003" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:28.79" heatid="27005" lane="3" />
                <ENTRY eventid="39" entrytime="00:00:27.64" heatid="39004" lane="3" />
                <ENTRY eventid="14" entrytime="00:01:06.45" heatid="14001" lane="6" />
                <ENTRY eventid="32" entrytime="00:01:00.57" heatid="32001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="492" eventid="1" swimtime="00:01:06.45" lane="3" heatid="1004" points="572" />
                <RESULT resultid="493" eventid="11" swimtime="00:01:00.57" lane="4" heatid="11003" points="622" />
                <RESULT resultid="816" eventid="14" swimtime="00:01:03.78" lane="6" heatid="14001" points="647" />
                <RESULT resultid="494" eventid="27" swimtime="00:00:29.19" lane="3" heatid="27005" points="586" />
                <RESULT resultid="868" eventid="32" swimtime="00:01:02.23" lane="2" heatid="32001" points="573" />
                <RESULT resultid="495" eventid="39" swimtime="00:00:28.00" lane="3" heatid="39004" points="599" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="2013-01-01" gender="M" lastname="Hanf" firstname="Leandro" license="464263" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:48.25" heatid="4002" lane="1" />
                <ENTRY eventid="12" entrytime="00:01:16.72" heatid="12001" lane="7" />
                <ENTRY eventid="24" entrytime="00:03:09.22" heatid="24001" lane="7" />
                <ENTRY eventid="28" entrytime="00:00:40.16" heatid="28001" lane="4" />
                <ENTRY eventid="36" entrytime="00:01:20.78" heatid="36001" lane="5" />
                <ENTRY eventid="44" entrytime="00:00:48.90" heatid="44001" lane="3" />
                <ENTRY eventid="46" entrytime="00:05:45.18" heatid="46001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="496" eventid="4" swimtime="00:02:40.99" lane="1" heatid="4002" points="254">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="497" eventid="12" swimtime="00:01:12.69" lane="7" heatid="12001" points="260" />
                <RESULT resultid="498" eventid="24" swimtime="00:03:01.66" lane="7" heatid="24001" points="247">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="499" eventid="28" swimtime="00:00:39.23" lane="4" heatid="28001" points="182" />
                <RESULT resultid="500" eventid="36" swimtime="00:01:19.29" lane="5" heatid="36001" points="275" />
                <RESULT resultid="501" eventid="44" swimtime="00:00:45.53" lane="3" heatid="44001" points="185" />
                <RESULT resultid="502" eventid="46" swimtime="00:05:37.54" lane="5" heatid="46001" points="277">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.10" />
                    <SPLIT distance="200" swimtime="00:02:47.10" />
                    <SPLIT distance="300" swimtime="00:04:14.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2009-01-01" gender="F" lastname="Karpa" firstname="Leonor" license="399381" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:07.74" heatid="1004" lane="6" />
                <ENTRY eventid="11" entrytime="00:01:01.72" heatid="11005" lane="2" />
                <ENTRY eventid="27" entrytime="00:00:29.99" heatid="27005" lane="8" />
                <ENTRY eventid="39" entrytime="00:00:28.41" heatid="39004" lane="8" />
                <ENTRY eventid="14" entrytime="00:01:08.78" heatid="14000" lane="0" />
                <ENTRY eventid="32" entrytime="00:01:02.40" heatid="32001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="503" eventid="1" swimtime="00:01:08.78" lane="6" heatid="1004" points="516" />
                <RESULT resultid="504" eventid="11" swimtime="00:01:02.40" lane="2" heatid="11005" points="569" />
                <RESULT resultid="811" eventid="14" status="WDR" swimtime="00:00:00.00" lane="0" heatid="14000" />
                <RESULT resultid="505" eventid="27" swimtime="00:00:30.30" lane="8" heatid="27005" points="524" />
                <RESULT resultid="869" eventid="32" swimtime="00:01:03.14" lane="7" heatid="32001" points="549" />
                <RESULT resultid="506" eventid="39" swimtime="00:00:28.68" lane="8" heatid="39004" points="557" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="2013-01-01" gender="F" lastname="Schröter" firstname="Lucia Sophie" license="440281" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:30.42" heatid="1001" lane="7" />
                <ENTRY eventid="7" entrytime="00:03:11.43" heatid="7001" lane="2" />
                <ENTRY eventid="21" entrytime="00:00:42.27" heatid="21001" lane="6" />
                <ENTRY eventid="23" entrytime="00:03:04.80" heatid="23001" lane="1" />
                <ENTRY eventid="35" entrytime="00:01:34.42" heatid="35001" lane="3" />
                <ENTRY eventid="45" entrytime="00:05:43.37" heatid="45002" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="507" eventid="1" swimtime="00:01:29.04" lane="7" heatid="1001" points="238" />
                <RESULT resultid="508" eventid="7" swimtime="00:03:02.45" lane="2" heatid="7001" points="307">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="509" eventid="21" swimtime="00:00:40.31" lane="6" heatid="21001" points="295" />
                <RESULT resultid="510" eventid="23" swimtime="00:03:00.69" lane="1" heatid="23001" points="340">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="511" eventid="35" swimtime="00:01:25.85" lane="3" heatid="35001" points="294" />
                <RESULT resultid="512" eventid="45" swimtime="00:05:36.89" lane="8" heatid="45002" points="341">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="200" swimtime="00:02:44.60" />
                    <SPLIT distance="300" swimtime="00:04:12.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110" birthdate="2008-01-01" gender="F" lastname="Weiß" firstname="Matilda" license="391730" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:09.76" heatid="3003" lane="6" />
                <ENTRY eventid="23" entrytime="00:02:31.15" heatid="23004" lane="4" />
                <ENTRY eventid="39" entrytime="00:00:28.69" heatid="39003" lane="3" />
                <ENTRY eventid="43" entrytime="00:00:39.88" heatid="43002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="513" eventid="3" swimtime="00:02:10.81" lane="6" heatid="3003" points="631">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="514" eventid="23" swimtime="00:02:33.53" lane="4" heatid="23004" points="554">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="515" eventid="39" swimtime="00:00:29.07" lane="3" heatid="39003" points="535" />
                <RESULT resultid="516" eventid="43" swimtime="00:00:41.12" lane="2" heatid="43002" points="356" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111" birthdate="2007-01-01" gender="M" lastname="Jonas" firstname="Melvin" license="405616" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:00.07" heatid="4004" lane="6" />
                <ENTRY eventid="12" entrytime="00:00:56.39" heatid="12003" lane="6" />
                <ENTRY eventid="46" entrytime="00:04:12.88" heatid="46003" lane="3" />
                <ENTRY eventid="34" entrytime="00:00:56.05" heatid="34001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="517" eventid="4" swimtime="00:01:59.22" lane="6" heatid="4004" points="626">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="518" eventid="12" swimtime="00:00:56.05" lane="6" heatid="12003" points="567" />
                <RESULT resultid="887" eventid="34" swimtime="00:00:56.43" lane="8" heatid="34001" points="555" />
                <RESULT resultid="519" eventid="46" swimtime="00:04:13.43" lane="3" heatid="46003" points="654">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.63" />
                    <SPLIT distance="200" swimtime="00:02:04.17" />
                    <SPLIT distance="300" swimtime="00:03:09.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="112" birthdate="2011-01-01" gender="F" lastname="Rockstroh" firstname="Mira Lysann" license="420406" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:13.51" heatid="3003" lane="8" />
                <ENTRY eventid="11" entrytime="00:01:02.33" heatid="11004" lane="2" />
                <ENTRY eventid="21" entrytime="00:00:33.74" heatid="21002" lane="4" />
                <ENTRY eventid="39" entrytime="00:00:28.97" heatid="39003" lane="2" />
                <ENTRY eventid="43" entrytime="00:00:43.56" heatid="43001" lane="5" />
                <ENTRY eventid="31" entrytime="00:01:01.48" heatid="31001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="520" eventid="3" swimtime="00:02:14.02" lane="8" heatid="3003" points="587">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="521" eventid="11" swimtime="00:01:01.48" lane="2" heatid="11004" points="595" />
                <RESULT resultid="522" eventid="21" swimtime="00:00:33.99" lane="4" heatid="21002" points="493" />
                <RESULT resultid="860" eventid="31" swimtime="00:01:01.81" lane="2" heatid="31001" points="585" />
                <RESULT resultid="523" eventid="39" swimtime="00:00:28.83" lane="2" heatid="39003" points="549" />
                <RESULT resultid="524" eventid="43" swimtime="00:00:38.12" lane="5" heatid="43001" points="447" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113" birthdate="2013-01-01" gender="F" lastname="Müller" firstname="Nele" license="449563" nation="GER">
              <ENTRIES>
                <ENTRY eventid="3" entrytime="00:02:34.63" heatid="3001" lane="5" />
                <ENTRY eventid="11" entrytime="00:01:08.30" heatid="11002" lane="4" />
                <ENTRY eventid="21" entrytime="00:00:37.88" heatid="21002" lane="8" />
                <ENTRY eventid="23" entrytime="00:02:51.71" heatid="23001" lane="4" />
                <ENTRY eventid="27" entrytime="00:00:34.12" heatid="27002" lane="5" />
                <ENTRY eventid="35" entrytime="00:01:23.40" heatid="35002" lane="7" />
                <ENTRY eventid="45" entrytime="00:05:36.26" heatid="45002" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="525" eventid="3" swimtime="00:02:33.86" lane="5" heatid="3001" points="388">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="526" eventid="11" swimtime="00:01:08.20" lane="4" heatid="11002" points="435" />
                <RESULT resultid="527" eventid="21" swimtime="00:00:37.60" lane="8" heatid="21002" points="364" />
                <RESULT resultid="528" eventid="23" swimtime="00:02:51.40" lane="4" heatid="23001" points="398">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="529" eventid="27" swimtime="00:00:34.75" lane="5" heatid="27002" points="347" />
                <RESULT resultid="530" eventid="35" swimtime="00:01:21.95" lane="7" heatid="35002" points="338" />
                <RESULT resultid="531" eventid="45" swimtime="00:05:26.40" lane="7" heatid="45002" points="375">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.86" />
                    <SPLIT distance="200" swimtime="00:02:39.99" />
                    <SPLIT distance="300" swimtime="00:04:05.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="114" birthdate="2014-01-01" gender="M" lastname="Bredau" firstname="Nuri" license="470040" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:58.40" heatid="4001" lane="3" />
                <ENTRY eventid="12" entrytime="00:01:20.32" heatid="12001" lane="8" />
                <ENTRY eventid="22" entrytime="00:00:44.08" heatid="22001" lane="3" />
                <ENTRY eventid="24" entrytime="00:03:16.25" heatid="24001" lane="8" />
                <ENTRY eventid="28" entrytime="00:00:50.26" heatid="28001" lane="5" />
                <ENTRY eventid="36" entrytime="00:01:37.48" heatid="36001" lane="7" />
                <ENTRY eventid="46" entrytime="00:06:07.15" heatid="46001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="532" eventid="4" swimtime="00:02:46.37" lane="3" heatid="4001" points="230">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="533" eventid="12" swimtime="00:01:14.84" lane="8" heatid="12001" points="238" />
                <RESULT resultid="534" eventid="22" swimtime="00:00:42.19" lane="3" heatid="22001" points="173" />
                <RESULT resultid="535" eventid="24" swimtime="00:03:07.52" lane="8" heatid="24001" points="224">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="536" eventid="28" swimtime="00:00:39.14" lane="5" heatid="28001" points="184" />
                <RESULT resultid="537" eventid="36" swimtime="00:01:29.83" lane="7" heatid="36001" points="189" />
                <RESULT resultid="538" eventid="46" swimtime="00:05:57.68" lane="6" heatid="46001" points="232">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="200" swimtime="00:02:57.40" />
                    <SPLIT distance="300" swimtime="00:04:30.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="115" birthdate="2011-01-01" gender="M" lastname="Erhard" firstname="Ole" license="423576" nation="GER">
              <ENTRIES>
                <ENTRY eventid="12" entrytime="00:01:02.50" heatid="12002" lane="3" />
                <ENTRY eventid="24" entrytime="00:02:32.74" heatid="24002" lane="4" />
                <ENTRY eventid="36" entrytime="00:01:08.14" heatid="36004" lane="2" />
                <ENTRY eventid="49" entrytime="00:01:08.18" heatid="49001" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="539" eventid="12" swimtime="00:01:01.58" lane="3" heatid="12002" points="427" />
                <RESULT resultid="540" eventid="24" swimtime="00:02:35.71" lane="4" heatid="24002" points="392">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="541" eventid="36" swimtime="00:01:08.18" lane="2" heatid="36004" points="433" />
                <RESULT resultid="906" eventid="49" swimtime="00:01:07.98" lane="7" heatid="49001" points="437" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="116" birthdate="2013-01-01" gender="F" lastname="Gebhardt" firstname="Pauline" license="445340" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:42.81" heatid="5002" lane="7" />
                <ENTRY eventid="11" entrytime="00:01:03.98" heatid="11005" lane="1" />
                <ENTRY eventid="21" entrytime="00:00:32.81" heatid="21003" lane="8" />
                <ENTRY eventid="27" entrytime="00:00:31.86" heatid="27003" lane="3" />
                <ENTRY eventid="37" entrytime="00:03:00.00" heatid="37001" lane="4" />
                <ENTRY eventid="31" entrytime="00:01:03.71" heatid="31001" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="542" eventid="5" swimtime="00:01:25.73" lane="7" heatid="5002" points="418" />
                <RESULT resultid="543" eventid="11" swimtime="00:01:03.71" lane="1" heatid="11005" points="534" />
                <RESULT resultid="544" eventid="21" swimtime="00:00:33.66" lane="8" heatid="21003" points="508" />
                <RESULT resultid="545" eventid="27" swimtime="00:00:33.31" lane="3" heatid="27003" points="394" />
                <RESULT resultid="862" eventid="31" swimtime="00:01:06.97" lane="1" heatid="31001" points="460" />
                <RESULT resultid="546" eventid="37" status="WDR" swimtime="00:00:00.00" lane="4" heatid="37001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="117" birthdate="2012-01-01" gender="F" lastname="Köhler" firstname="Swenja" license="434391" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:33.81" heatid="5001" lane="2" />
                <ENTRY eventid="11" entrytime="00:01:12.60" heatid="11002" lane="3" />
                <ENTRY eventid="21" entrytime="00:00:36.68" heatid="21002" lane="7" />
                <ENTRY eventid="29" entrytime="00:03:25.10" heatid="29001" lane="5" />
                <ENTRY eventid="39" entrytime="00:00:33.08" heatid="39002" lane="1" />
                <ENTRY eventid="45" entrytime="00:05:28.93" heatid="45002" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="547" eventid="5" swimtime="00:01:27.40" lane="2" heatid="5001" points="395" />
                <RESULT resultid="548" eventid="11" swimtime="00:01:11.57" lane="3" heatid="11002" points="377" />
                <RESULT resultid="549" eventid="21" swimtime="00:00:36.19" lane="7" heatid="21002" points="408" />
                <RESULT resultid="550" eventid="29" swimtime="00:03:07.68" lane="5" heatid="29001" points="393">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="551" eventid="39" swimtime="00:00:32.28" lane="1" heatid="39002" points="391" />
                <RESULT resultid="552" eventid="45" swimtime="00:05:21.00" lane="2" heatid="45002" points="394">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.34" />
                    <SPLIT distance="200" swimtime="00:02:39.00" />
                    <SPLIT distance="300" swimtime="00:04:01.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118" birthdate="2011-01-01" gender="M" lastname="Karpa" firstname="Thorben" license="407287" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:08.88" heatid="2005" lane="1" />
                <ENTRY eventid="24" entrytime="00:02:34.30" heatid="24002" lane="5" />
                <ENTRY eventid="28" entrytime="00:00:30.40" heatid="28004" lane="6" />
                <ENTRY eventid="42" entrytime="00:05:31.78" heatid="42003" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="553" eventid="2" swimtime="00:01:06.85" lane="1" heatid="2005" points="404" />
                <RESULT resultid="554" eventid="24" swimtime="00:02:30.15" lane="5" heatid="24002" points="437">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="555" eventid="28" swimtime="00:00:29.98" lane="6" heatid="28004" points="409" />
                <RESULT resultid="556" eventid="42" swimtime="00:05:17.81" lane="1" heatid="42003" points="444">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.27" />
                    <SPLIT distance="200" swimtime="00:02:29.65" />
                    <SPLIT distance="300" swimtime="00:04:06.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="119" birthdate="2013-01-01" gender="M" lastname="Götze" firstname="Vincent" license="448825" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:46.91" heatid="4002" lane="7" />
                <ENTRY eventid="12" entrytime="00:01:14.93" heatid="12001" lane="2" />
                <ENTRY eventid="22" entrytime="00:00:38.39" heatid="22001" lane="5" />
                <ENTRY eventid="24" entrytime="00:02:57.84" heatid="24001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="557" eventid="4" swimtime="00:02:34.31" lane="7" heatid="4002" points="288">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="558" eventid="12" swimtime="00:01:10.17" lane="2" heatid="12001" points="289" />
                <RESULT resultid="559" eventid="22" swimtime="00:00:37.58" lane="5" heatid="22001" points="246" />
                <RESULT resultid="560" eventid="24" swimtime="00:02:55.58" lane="2" heatid="24001" points="273">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Weixdorf" nation="GER" region="12" code="3366">
          <ATHLETES>
            <ATHLETE athleteid="3" birthdate="2007-01-01" gender="M" lastname="Koenig" firstname="Gabriel" license="333012" nation="GER">
              <ENTRIES>
                <ENTRY eventid="4" entrytime="00:02:04.42" heatid="4003" lane="4" />
                <ENTRY eventid="12" entrytime="00:00:56.90" heatid="12003" lane="2" />
                <ENTRY eventid="28" entrytime="00:00:27.65" heatid="28006" lane="8" />
                <ENTRY eventid="40" entrytime="00:00:25.97" heatid="40005" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="8" eventid="4" swimtime="00:02:08.55" lane="4" heatid="4003" points="499">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="9" eventid="12" swimtime="00:00:57.87" lane="2" heatid="12003" points="515" />
                <RESULT resultid="10" eventid="28" swimtime="00:00:28.16" lane="8" heatid="28006" points="494" />
                <RESULT resultid="11" eventid="40" swimtime="00:00:26.58" lane="8" heatid="40005" points="486" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SVV Plauen" nation="GER" region="12" code="6253">
          <ATHLETES>
            <ATHLETE athleteid="89" birthdate="2011-01-01" gender="M" lastname="Schwanke" firstname="Tim" license="423421">
              <ENTRIES>
                <ENTRY eventid="6" entrytime="00:01:18.11" heatid="6002" lane="3" />
                <ENTRY eventid="12" entrytime="00:00:59.56" heatid="12005" lane="1" />
                <ENTRY eventid="40" entrytime="00:00:26.89" heatid="40004" lane="2" />
                <ENTRY eventid="44" entrytime="00:00:34.58" heatid="44002" lane="4" />
                <ENTRY eventid="19" entrytime="00:01:15.45" heatid="19001" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="430" eventid="6" swimtime="00:01:15.45" lane="3" heatid="6002" points="428" />
                <RESULT resultid="431" eventid="12" swimtime="00:00:59.96" lane="1" heatid="12005" points="463" />
                <RESULT resultid="848" eventid="19" swimtime="00:01:16.75" lane="6" heatid="19001" points="407" />
                <RESULT resultid="432" eventid="40" swimtime="00:00:26.82" lane="2" heatid="40004" points="473" />
                <RESULT resultid="433" eventid="44" swimtime="00:00:34.79" lane="4" heatid="44002" points="415" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SWV TuR Dresden" nation="GER" region="12" code="3358">
          <ATHLETES>
            <ATHLETE athleteid="48" birthdate="2012-01-01" gender="M" lastname="Fischer" firstname="Lennox" license="445086" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:09:46.84" heatid="10002" lane="1" />
                <ENTRY eventid="22" entrytime="00:00:35.19" heatid="22002" lane="3" />
                <ENTRY eventid="28" entrytime="00:00:34.12" heatid="28003" lane="1" />
                <ENTRY eventid="46" entrytime="00:04:46.55" heatid="46002" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="238" eventid="10" swimtime="00:10:17.66" lane="1" heatid="10002" points="392">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.02" />
                    <SPLIT distance="200" swimtime="00:02:26.53" />
                    <SPLIT distance="300" swimtime="00:03:44.02" />
                    <SPLIT distance="400" swimtime="00:05:01.97" />
                    <SPLIT distance="500" swimtime="00:06:20.84" />
                    <SPLIT distance="600" swimtime="00:07:39.73" />
                    <SPLIT distance="700" swimtime="00:08:58.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="239" eventid="22" swimtime="00:00:35.26" lane="3" heatid="22002" points="297" />
                <RESULT resultid="240" eventid="28" swimtime="00:00:35.75" lane="1" heatid="28003" points="241" />
                <RESULT resultid="241" eventid="46" swimtime="00:04:56.64" lane="3" heatid="46002" points="408">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.73" />
                    <SPLIT distance="200" swimtime="00:02:24.17" />
                    <SPLIT distance="300" swimtime="00:03:40.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="USV TU Dresden e.V." nation="GER" region="12" code="3410">
          <ATHLETES>
            <ATHLETE athleteid="9" birthdate="2008-01-01" gender="F" lastname="Grammlich" firstname="Katharina" license="380800" nation="GER">
              <ENTRIES>
                <ENTRY eventid="5" entrytime="00:01:18.24" heatid="5003" lane="6" />
                <ENTRY eventid="21" entrytime="00:00:30.59" heatid="21003" lane="5" />
                <ENTRY eventid="35" entrytime="00:01:07.13" heatid="35003" lane="4" />
                <ENTRY eventid="43" entrytime="00:00:34.85" heatid="43003" lane="3" />
                <ENTRY eventid="18" entrytime="00:01:20.50" heatid="18001" lane="6" />
                <ENTRY eventid="48" entrytime="00:01:10.81" heatid="48001" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="35" eventid="5" swimtime="00:01:20.50" lane="6" heatid="5003" points="505" />
                <RESULT resultid="844" eventid="18" swimtime="00:01:19.65" lane="6" heatid="18001" points="521" />
                <RESULT resultid="36" eventid="21" swimtime="00:00:33.02" lane="5" heatid="21003" points="538" />
                <RESULT resultid="37" eventid="35" swimtime="00:01:10.81" lane="4" heatid="35003" points="525" />
                <RESULT resultid="38" eventid="43" swimtime="00:00:36.01" lane="3" heatid="43003" points="530" />
                <RESULT resultid="900" eventid="48" swimtime="00:01:12.28" lane="2" heatid="48001" points="493" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="10" birthdate="2012-01-01" gender="M" lastname="Kurlykov" firstname="Kirill" license="437629" nation="GER">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:10:41.30" heatid="10001" lane="6" />
                <ENTRY eventid="24" entrytime="00:02:38.32" heatid="24002" lane="6" />
                <ENTRY eventid="28" entrytime="00:00:32.54" heatid="28003" lane="4" />
                <ENTRY eventid="40" entrytime="00:00:29.90" heatid="40003" lane="8" />
                <ENTRY eventid="46" entrytime="00:05:24.60" heatid="46001" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="39" eventid="10" swimtime="00:10:28.82" lane="6" heatid="10001" points="371">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="200" swimtime="00:02:29.53" />
                    <SPLIT distance="300" swimtime="00:03:49.07" />
                    <SPLIT distance="400" swimtime="00:05:10.42" />
                    <SPLIT distance="500" swimtime="00:06:31.60" />
                    <SPLIT distance="600" swimtime="00:07:51.89" />
                    <SPLIT distance="700" swimtime="00:09:12.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="40" eventid="24" swimtime="00:02:41.09" lane="6" heatid="24002" points="354">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="41" eventid="28" swimtime="00:00:32.37" lane="4" heatid="28003" points="325" />
                <RESULT resultid="42" eventid="40" swimtime="00:00:29.99" lane="8" heatid="40003" points="338" />
                <RESULT resultid="43" eventid="46" swimtime="00:05:07.04" lane="4" heatid="46001" points="368">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.58" />
                    <SPLIT distance="200" swimtime="00:02:32.51" />
                    <SPLIT distance="300" swimtime="00:03:51.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="11" birthdate="2011-01-01" gender="M" lastname="Langner" firstname="Lukas" license="426678" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:13.06" heatid="2005" lane="8" />
                <ENTRY eventid="24" entrytime="00:02:28.27" heatid="24003" lane="6" />
                <ENTRY eventid="28" entrytime="00:00:31.20" heatid="28004" lane="8" />
                <ENTRY eventid="36" entrytime="00:01:07.93" heatid="36002" lane="6" />
                <ENTRY eventid="40" entrytime="00:00:28.59" heatid="40003" lane="6" />
                <ENTRY eventid="49" entrytime="00:01:10.56" heatid="49001" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="44" eventid="2" swimtime="00:01:07.28" lane="8" heatid="2005" points="397" />
                <RESULT resultid="45" eventid="24" swimtime="00:02:31.10" lane="6" heatid="24003" points="429">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="46" eventid="28" swimtime="00:00:30.59" lane="8" heatid="28004" points="385" />
                <RESULT resultid="47" eventid="36" swimtime="00:01:10.56" lane="6" heatid="36002" points="391" />
                <RESULT resultid="48" eventid="40" swimtime="00:00:28.57" lane="6" heatid="40003" points="392" />
                <RESULT resultid="908" eventid="49" swimtime="00:01:08.77" lane="8" heatid="49001" points="422" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="12" birthdate="2012-01-01" gender="F" lastname="Dittel" firstname="Magdalena" license="437623" nation="GER">
              <ENTRIES>
                <ENTRY eventid="1" entrytime="00:01:13.77" heatid="1002" lane="1" />
                <ENTRY eventid="11" entrytime="00:01:02.61" heatid="11003" lane="2" />
                <ENTRY eventid="21" entrytime="00:00:32.16" heatid="21003" lane="7" />
                <ENTRY eventid="35" entrytime="00:01:09.61" heatid="35003" lane="3" />
                <ENTRY eventid="39" entrytime="00:00:29.70" heatid="39002" lane="4" />
                <ENTRY eventid="47" entrytime="00:01:09.45" heatid="47001" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="49" eventid="1" swimtime="00:01:14.19" lane="1" heatid="1002" points="411" />
                <RESULT resultid="50" eventid="11" swimtime="00:01:04.43" lane="2" heatid="11003" points="516" />
                <RESULT resultid="51" eventid="21" swimtime="00:00:32.48" lane="7" heatid="21003" points="565" />
                <RESULT resultid="52" eventid="35" swimtime="00:01:09.45" lane="3" heatid="35003" points="556" />
                <RESULT resultid="53" eventid="39" swimtime="00:00:29.93" lane="4" heatid="39002" points="490" />
                <RESULT resultid="889" eventid="47" swimtime="00:01:10.70" lane="5" heatid="47001" points="527" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="W98 Hannover" nation="GER" region="9" code="6661">
          <ATHLETES>
            <ATHLETE athleteid="64" birthdate="2014-01-01" gender="M" lastname="Müller" firstname="Jannis" license="465820" nation="GER">
              <ENTRIES>
                <ENTRY eventid="2" entrytime="00:01:18.48" heatid="2003" lane="8" />
                <ENTRY eventid="12" entrytime="00:01:07.05" heatid="12002" lane="2" />
                <ENTRY eventid="26" entrytime="00:20:00.00" heatid="26002" lane="3" />
                <ENTRY eventid="42" entrytime="00:05:59.44" heatid="42002" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT resultid="306" eventid="2" swimtime="00:01:18.50" lane="8" heatid="2003" points="249" />
                <RESULT resultid="307" eventid="12" swimtime="00:01:05.53" lane="2" heatid="12002" points="355" />
                <RESULT resultid="308" eventid="26" swimtime="00:19:37.35" lane="3" heatid="26002" points="404">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="200" swimtime="00:02:25.80" />
                    <SPLIT distance="300" swimtime="00:03:43.92" />
                    <SPLIT distance="400" swimtime="00:05:02.71" />
                    <SPLIT distance="500" swimtime="00:06:23.05" />
                    <SPLIT distance="600" swimtime="00:07:42.15" />
                    <SPLIT distance="700" swimtime="00:09:01.52" />
                    <SPLIT distance="800" swimtime="00:10:21.01" />
                    <SPLIT distance="900" swimtime="00:11:41.08" />
                    <SPLIT distance="1000" swimtime="00:13:00.95" />
                    <SPLIT distance="1100" swimtime="00:14:20.14" />
                    <SPLIT distance="1200" swimtime="00:15:40.03" />
                    <SPLIT distance="1300" swimtime="00:17:00.17" />
                    <SPLIT distance="1400" swimtime="00:18:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="309" eventid="42" swimtime="00:05:54.12" lane="5" heatid="42002" points="321">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.54" />
                    <SPLIT distance="200" swimtime="00:02:51.59" />
                    <SPLIT distance="300" swimtime="00:04:35.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
