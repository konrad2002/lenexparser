﻿<?xml version="1.0" encoding="UTF-8"?>
<LENEX revisiondate="2024-12-02" created="2025-12-17T06:29:01" version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Dresdner SC 1898" version="11.83082">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Dresden" name="33. Internationales Dresdner Christstollen-Schwimmfest" course="LCM" deadline="2025-12-08" hostclub="Dresdner SC 1898" hostclub.url="https://schwimmen.dsc1898.de/" organizer="Dresdner SC 1898" organizer.url="https://schwimmen.dsc1898.de/" result.url="https://live.swimrankings.net/45267/" startmethod="1" status="SEEDED" timing="AUTOMATIC" touchpad="BOTHSIDE" masters="F" state="SN" nation="GER" hytek.courseorder="L">
      <AGEDATE value="2025-01-01" type="YEAR" />
      <POOL name="SSK Freiberger Platz" lanemin="1" lanemax="8" />
      <FACILITY city="Dresden" name="SSK Freiberger Platz" nation="GER" state="SN" />
      <POINTTABLE pointtableid="3018" name="AQUA Point Scoring" version="2025" />
      <QUALIFY from="2025-01-01" until="2025-12-09" conversion="NON_CONFORMING_LAST" />
      <CONTACT city="Dresden" email="meldung.schwimmen@dsc1898.de" name="Silke Rößler" street="Magdeburger Straße 12" zip="01067" />
      <SESSIONS>
        <SESSION date="2025-12-19" daytime="15:30" endtime="21:53" number="1" officialmeeting="15:00" status="SEEDED" warmupfrom="14:30">
          <EVENTS>
            <EVENT eventid="1063" daytime="15:30" gender="F" number="1" order="1" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1065" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1066" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1067" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1068" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1069" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1070" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1071" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1072" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="39994" daytime="15:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="39995" daytime="15:37" number="2" order="2" status="SEEDED" />
                <HEAT heatid="39996" daytime="15:43" number="3" order="3" status="SEEDED" />
                <HEAT heatid="39997" daytime="15:50" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1073" daytime="15:56" gender="M" number="2" order="2" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1074" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1075" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1076" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1077" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1078" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1079" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1080" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1081" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1082" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="39998" daytime="15:56" number="1" order="1" status="SEEDED" />
                <HEAT heatid="39999" daytime="16:03" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40000" daytime="16:10" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40001" daytime="16:16" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40002" daytime="16:22" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1083" daytime="16:27" gender="F" number="3" order="3" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1085" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1086" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1087" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1088" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1089" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1090" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1091" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1092" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40003" daytime="16:27" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40004" daytime="16:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40005" daytime="16:53" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40006" daytime="17:05" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40007" daytime="17:17" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40008" daytime="17:28" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40009" daytime="17:40" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40010" daytime="17:51" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40011" daytime="18:02" number="9" order="9" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1093" daytime="18:12" gender="M" number="4" order="4" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1094" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1095" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1096" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1097" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1098" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1099" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1100" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1101" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1102" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40012" daytime="18:12" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40013" daytime="18:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40014" daytime="18:38" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40015" daytime="18:49" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40016" daytime="19:00" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40017" daytime="19:11" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40018" daytime="19:22" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40019" daytime="19:32" number="8" order="8" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1103" daytime="19:42" gender="F" number="5" order="5" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1105" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1106" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1107" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1108" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1109" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1110" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1111" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1112" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40020" daytime="19:42" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40021" daytime="20:04" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1113" daytime="20:27" gender="M" number="6" order="6" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1115" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1116" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1117" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1118" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1119" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1120" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1121" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1122" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40022" daytime="20:27" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40023" daytime="20:50" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40024" daytime="21:12" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40025" daytime="21:33" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="55" />
            <JUDGE officialid="85" />
            <JUDGE officialid="62" />
            <JUDGE officialid="69" />
            <JUDGE officialid="12" />
            <JUDGE officialid="78" />
            <JUDGE officialid="35999" />
            <JUDGE officialid="36003" />
            <JUDGE officialid="52" />
            <JUDGE officialid="36007" />
            <JUDGE officialid="25" />
            <JUDGE officialid="36004" />
            <JUDGE officialid="14" />
            <JUDGE officialid="20596" />
            <JUDGE officialid="36006" />
            <JUDGE officialid="35861" />
            <JUDGE officialid="20598" />
            <JUDGE officialid="70" />
            <JUDGE officialid="16" />
            <JUDGE officialid="36001" />
            <JUDGE officialid="35865" />
            <JUDGE officialid="20599" />
            <JUDGE officialid="79" />
            <JUDGE officialid="36000" />
            <JUDGE officialid="36000" />
            <JUDGE officialid="36005" />
            <JUDGE officialid="36005" />
            <JUDGE officialid="36002" />
            <JUDGE officialid="36002" />
            <JUDGE officialid="20597" />
            <JUDGE officialid="20597" />
          </JUDGES>
        </SESSION>
        <SESSION date="2025-12-20" daytime="09:30" endtime="13:54" number="2" officialmeeting="09:00" status="SEEDED" warmupfrom="08:30">
          <EVENTS>
            <EVENT eventid="1123" daytime="09:30" gender="F" number="7" order="1" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1124" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1125" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1126" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1127" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1128" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1129" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1130" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1131" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1132" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40026" daytime="09:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40027" daytime="09:31" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40028" daytime="09:32" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40029" daytime="09:33" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40030" daytime="09:35" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40031" daytime="09:36" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40032" daytime="09:37" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40033" daytime="09:38" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40034" daytime="09:39" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40035" daytime="09:40" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40036" daytime="09:41" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40037" daytime="09:42" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40038" daytime="09:43" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40039" daytime="09:44" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40040" daytime="09:45" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40041" daytime="09:46" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40042" daytime="09:47" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40043" daytime="09:48" number="18" order="18" status="SEEDED" />
                <HEAT heatid="40044" daytime="09:49" number="19" order="19" status="SEEDED" />
                <HEAT heatid="40045" daytime="09:50" number="20" order="20" status="SEEDED" />
                <HEAT heatid="40046" daytime="09:51" number="21" order="21" status="SEEDED" />
                <HEAT heatid="40047" daytime="09:52" number="22" order="22" status="SEEDED" />
                <HEAT heatid="40048" daytime="09:53" number="23" order="23" status="SEEDED" />
                <HEAT heatid="40049" daytime="09:54" number="24" order="24" status="SEEDED" />
                <HEAT heatid="40050" daytime="09:55" number="25" order="25" status="SEEDED" />
                <HEAT heatid="40051" daytime="09:56" number="26" order="26" status="SEEDED" />
                <HEAT heatid="40052" daytime="09:57" number="27" order="27" status="SEEDED" />
                <HEAT heatid="40053" daytime="09:58" number="28" order="28" status="SEEDED" />
                <HEAT heatid="40054" daytime="09:59" number="29" order="29" status="SEEDED" />
                <HEAT heatid="40055" daytime="10:00" number="30" order="30" status="SEEDED" />
                <HEAT heatid="40056" daytime="10:01" number="31" order="31" status="SEEDED" />
                <HEAT heatid="40057" daytime="10:02" number="32" order="32" status="SEEDED" />
                <HEAT heatid="40058" daytime="10:03" number="33" order="33" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1133" daytime="10:04" gender="M" number="8" order="2" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1134" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1135" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1136" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1137" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1138" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1139" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1140" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1141" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1142" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40059" daytime="10:04" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40060" daytime="10:06" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40061" daytime="10:07" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40062" daytime="10:08" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40063" daytime="10:09" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40064" daytime="10:10" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40065" daytime="10:11" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40066" daytime="10:12" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40067" daytime="10:13" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40068" daytime="10:14" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40069" daytime="10:15" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40070" daytime="10:16" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40071" daytime="10:17" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40072" daytime="10:18" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40073" daytime="10:19" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40074" daytime="10:20" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40075" daytime="10:21" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40076" daytime="10:22" number="18" order="18" status="SEEDED" />
                <HEAT heatid="40077" daytime="10:23" number="19" order="19" status="SEEDED" />
                <HEAT heatid="40078" daytime="10:24" number="20" order="20" status="SEEDED" />
                <HEAT heatid="40079" daytime="10:25" number="21" order="21" status="SEEDED" />
                <HEAT heatid="40080" daytime="10:26" number="22" order="22" status="SEEDED" />
                <HEAT heatid="40081" daytime="10:27" number="23" order="23" status="SEEDED" />
                <HEAT heatid="40082" daytime="10:28" number="24" order="24" status="SEEDED" />
                <HEAT heatid="40083" daytime="10:29" number="25" order="25" status="SEEDED" />
                <HEAT heatid="40084" daytime="10:30" number="26" order="26" status="SEEDED" />
                <HEAT heatid="40085" daytime="10:31" number="27" order="27" status="SEEDED" />
                <HEAT heatid="40086" daytime="10:32" number="28" order="28" status="SEEDED" />
                <HEAT heatid="40087" daytime="10:33" number="29" order="29" status="SEEDED" />
                <HEAT heatid="40088" daytime="10:34" number="30" order="30" status="SEEDED" />
                <HEAT heatid="40089" daytime="10:35" number="31" order="31" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1143" daytime="10:36" gender="F" number="9" order="3" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1144" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1145" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1146" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1147" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1148" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1149" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1150" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1151" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1152" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40090" daytime="10:36" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40091" daytime="10:42" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40092" daytime="10:46" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40093" daytime="10:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40094" daytime="10:54" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40095" daytime="10:58" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40096" daytime="11:01" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40097" daytime="11:05" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40098" daytime="11:09" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40099" daytime="11:12" number="10" order="10" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1153" daytime="11:16" gender="M" number="10" order="4" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1154" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1155" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1156" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1157" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1158" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1159" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1160" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1161" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1162" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40101" daytime="11:16" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40102" daytime="11:20" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40103" daytime="11:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40104" daytime="11:29" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40105" daytime="11:32" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40106" daytime="11:36" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40107" daytime="11:40" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40108" daytime="11:43" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40109" daytime="11:47" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40110" daytime="11:50" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40111" daytime="11:53" number="11" order="11" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1163" daytime="11:56" gender="F" number="11" order="5" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1164" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1165" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1166" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1167" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1168" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1169" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1170" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1171" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1172" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40112" daytime="11:56" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40113" daytime="12:01" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40114" daytime="12:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40115" daytime="12:08" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40116" daytime="12:12" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40117" daytime="12:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40118" daytime="12:19" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40119" daytime="12:22" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40120" daytime="12:26" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40121" daytime="12:29" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40122" daytime="12:32" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40123" daytime="12:36" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40124" daytime="12:39" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40125" daytime="12:42" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40126" daytime="12:45" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40127" daytime="12:48" number="16" order="16" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1173" daytime="12:51" gender="M" number="12" order="6" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1174" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1175" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1176" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1177" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1178" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1179" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1180" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1181" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1182" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40128" daytime="12:51" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40129" daytime="12:55" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40130" daytime="12:59" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40131" daytime="13:03" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40132" daytime="13:06" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40133" daytime="13:10" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40134" daytime="13:13" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40135" daytime="13:17" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40136" daytime="13:20" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40137" daytime="13:23" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40138" daytime="13:26" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40139" daytime="13:30" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40140" daytime="13:33" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40141" daytime="13:35" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40142" daytime="13:38" number="15" order="15" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1183" daytime="13:41" gender="F" number="13" order="7" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE value="900" />
              <HEATS>
                <HEAT heatid="40143" daytime="13:41" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40144" daytime="13:44" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1185" daytime="13:48" gender="M" number="14" order="8" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE value="900" />
              <HEATS>
                <HEAT heatid="40145" daytime="13:48" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40146" daytime="13:51" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="55" />
            <JUDGE officialid="85" />
            <JUDGE officialid="62" />
            <JUDGE officialid="69" />
            <JUDGE officialid="12" />
            <JUDGE officialid="78" />
            <JUDGE officialid="16" />
            <JUDGE officialid="36002" />
            <JUDGE officialid="52" />
            <JUDGE officialid="36007" />
            <JUDGE officialid="25" />
            <JUDGE officialid="36003" />
            <JUDGE officialid="13" />
            <JUDGE officialid="20596" />
            <JUDGE officialid="35999" />
            <JUDGE officialid="36000" />
            <JUDGE officialid="20598" />
            <JUDGE officialid="20599" />
            <JUDGE officialid="35863" />
            <JUDGE officialid="35861" />
            <JUDGE officialid="70" />
            <JUDGE officialid="20597" />
            <JUDGE officialid="79" />
            <JUDGE officialid="36001" />
            <JUDGE officialid="36001" />
            <JUDGE officialid="36004" />
            <JUDGE officialid="36004" />
            <JUDGE officialid="35861" />
            <JUDGE officialid="35861" />
            <JUDGE officialid="14" />
            <JUDGE officialid="14" />
          </JUDGES>
        </SESSION>
        <SESSION date="2025-12-20" daytime="14:25" endtime="19:43" number="3" status="SEEDED">
          <EVENTS>
            <EVENT eventid="1187" daytime="14:25" gender="F" number="15" order="1" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1188" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1189" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1190" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1191" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1192" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1193" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1194" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1195" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1196" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40147" daytime="14:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40148" daytime="14:29" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40149" daytime="14:32" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40150" daytime="14:36" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1197" daytime="14:39" gender="M" number="16" order="2" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1198" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1199" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1200" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1201" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1202" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1203" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1204" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1205" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1206" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40151" daytime="14:39" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40152" daytime="14:43" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40153" daytime="14:47" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40154" daytime="14:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40155" daytime="14:53" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40156" daytime="14:56" number="6" order="6" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1207" daytime="14:59" gender="F" number="17" order="3" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1208" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1209" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1210" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1211" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1212" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1213" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1214" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1215" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1216" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40157" daytime="14:59" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40158" daytime="15:01" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40159" daytime="15:02" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40160" daytime="15:03" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40161" daytime="15:04" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40162" daytime="15:06" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40163" daytime="15:07" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40164" daytime="15:08" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40165" daytime="15:09" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40166" daytime="15:10" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40167" daytime="15:12" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40168" daytime="15:13" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40169" daytime="15:14" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40170" daytime="15:15" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40171" daytime="15:16" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40172" daytime="15:17" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40173" daytime="15:19" number="17" order="17" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1217" daytime="15:20" gender="M" number="18" order="4" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1218" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1219" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1220" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1221" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1222" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1223" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1224" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1225" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1226" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40174" daytime="15:20" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40175" daytime="15:21" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40176" daytime="15:23" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40177" daytime="15:24" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40178" daytime="15:25" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40179" daytime="15:26" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40180" daytime="15:28" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40181" daytime="15:29" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40182" daytime="15:30" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40183" daytime="15:31" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40184" daytime="15:32" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40185" daytime="15:33" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40186" daytime="15:34" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40187" daytime="15:35" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40188" daytime="15:36" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40189" daytime="15:37" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40190" daytime="15:38" number="17" order="17" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1227" daytime="15:40" gender="F" number="19" order="5" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1228" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1229" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1230" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1231" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1232" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1233" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1234" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1235" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1236" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40191" daytime="15:40" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40192" daytime="15:42" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40193" daytime="15:44" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40194" daytime="15:46" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40195" daytime="15:48" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40196" daytime="15:50" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40197" daytime="15:52" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40198" daytime="15:54" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40199" daytime="15:56" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40200" daytime="15:58" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40201" daytime="16:00" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40202" daytime="16:02" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40203" daytime="16:04" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40204" daytime="16:05" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40205" daytime="16:07" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40206" daytime="16:09" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40207" daytime="16:11" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40208" daytime="16:13" number="18" order="18" status="SEEDED" />
                <HEAT heatid="40209" daytime="16:14" number="19" order="19" status="SEEDED" />
                <HEAT heatid="40210" daytime="16:16" number="20" order="20" status="SEEDED" />
                <HEAT heatid="40211" daytime="16:18" number="21" order="21" status="SEEDED" />
                <HEAT heatid="40212" daytime="16:20" number="22" order="22" status="SEEDED" />
                <HEAT heatid="40213" daytime="16:21" number="23" order="23" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1237" daytime="16:23" gender="M" number="20" order="6" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1238" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1239" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1240" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1241" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1242" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1243" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1244" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1245" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1246" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40214" daytime="16:23" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40215" daytime="16:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40216" daytime="16:28" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40217" daytime="16:30" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40218" daytime="16:32" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40219" daytime="16:34" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40220" daytime="16:35" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40221" daytime="16:37" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40222" daytime="16:39" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40223" daytime="16:41" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40224" daytime="16:43" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40225" daytime="16:45" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40226" daytime="16:46" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40227" daytime="16:48" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40228" daytime="16:50" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40229" daytime="16:52" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40230" daytime="16:53" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40231" daytime="16:55" number="18" order="18" status="SEEDED" />
                <HEAT heatid="40232" daytime="16:57" number="19" order="19" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1247" daytime="16:58" gender="F" number="21" order="7" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1248" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1249" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1250" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1251" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1252" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1253" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1254" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1255" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1256" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40233" daytime="16:58" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40234" daytime="17:06" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40235" daytime="17:13" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40236" daytime="17:19" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40237" daytime="17:26" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40238" daytime="17:32" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40239" daytime="17:38" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40240" daytime="17:44" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40241" daytime="17:49" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40242" daytime="17:55" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40243" daytime="18:01" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40244" daytime="18:06" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40245" daytime="18:12" number="13" order="13" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1257" daytime="18:17" gender="M" number="22" order="8" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1258" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1259" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1260" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1261" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1262" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1263" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1264" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1265" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1266" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40246" daytime="18:17" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40247" daytime="18:24" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40248" daytime="18:31" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40249" daytime="18:37" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40250" daytime="18:43" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40251" daytime="18:49" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40252" daytime="18:55" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40253" daytime="19:01" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40254" daytime="19:07" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40255" daytime="19:12" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40256" daytime="19:18" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40257" daytime="19:23" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40258" daytime="19:28" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40259" daytime="19:33" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40260" daytime="19:38" number="15" order="15" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2025-12-21" daytime="09:00" endtime="13:36" number="4" officialmeeting="08:30" status="SEEDED" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1267" daytime="09:00" gender="F" number="23" order="1" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1268" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1269" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1270" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1271" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1272" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1273" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1274" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1275" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1276" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40261" daytime="09:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40262" daytime="09:02" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40263" daytime="09:04" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40264" daytime="09:06" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40265" daytime="09:08" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40266" daytime="09:09" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40267" daytime="09:11" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40268" daytime="09:13" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40269" daytime="09:15" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40270" daytime="09:16" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40271" daytime="09:18" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40272" daytime="09:20" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40273" daytime="09:21" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40274" daytime="09:23" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40275" daytime="09:25" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40276" daytime="09:26" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40277" daytime="09:28" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40278" daytime="09:30" number="18" order="18" status="SEEDED" />
                <HEAT heatid="40279" daytime="09:31" number="19" order="19" status="SEEDED" />
                <HEAT heatid="40280" daytime="09:33" number="20" order="20" status="SEEDED" />
                <HEAT heatid="40281" daytime="09:35" number="21" order="21" status="SEEDED" />
                <HEAT heatid="40282" daytime="09:36" number="22" order="22" status="SEEDED" />
                <HEAT heatid="40283" daytime="09:38" number="23" order="23" status="SEEDED" />
                <HEAT heatid="40284" daytime="09:39" number="24" order="24" status="SEEDED" />
                <HEAT heatid="40285" daytime="09:41" number="25" order="25" status="SEEDED" />
                <HEAT heatid="40286" daytime="09:42" number="26" order="26" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1277" daytime="09:44" gender="M" number="24" order="2" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1278" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1279" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1280" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1281" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1282" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1283" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1284" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1285" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1286" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40287" daytime="09:44" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40288" daytime="09:46" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40289" daytime="09:48" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40290" daytime="09:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40291" daytime="09:52" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40292" daytime="09:54" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40293" daytime="09:55" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40294" daytime="09:57" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40295" daytime="09:59" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40296" daytime="10:01" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40297" daytime="10:02" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40298" daytime="10:04" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40299" daytime="10:06" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40300" daytime="10:07" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40301" daytime="10:09" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40302" daytime="10:10" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40303" daytime="10:12" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40304" daytime="10:13" number="18" order="18" status="SEEDED" />
                <HEAT heatid="40305" daytime="10:15" number="19" order="19" status="SEEDED" />
                <HEAT heatid="40306" daytime="10:16" number="20" order="20" status="SEEDED" />
                <HEAT heatid="40307" daytime="10:18" number="21" order="21" status="SEEDED" />
                <HEAT heatid="40308" daytime="10:19" number="22" order="22" status="SEEDED" />
                <HEAT heatid="40309" daytime="10:21" number="23" order="23" status="SEEDED" />
                <HEAT heatid="40310" daytime="10:22" number="24" order="24" status="SEEDED" />
                <HEAT heatid="40311" daytime="10:24" number="25" order="25" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1287" daytime="10:25" gender="F" number="25" order="3" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1288" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1289" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1290" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1291" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1292" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1293" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1294" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1295" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1296" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40312" daytime="10:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40313" daytime="10:27" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40314" daytime="10:28" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40315" daytime="10:29" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40316" daytime="10:30" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40317" daytime="10:31" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40318" daytime="10:32" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40319" daytime="10:33" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40320" daytime="10:34" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40321" daytime="10:35" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40322" daytime="10:37" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40323" daytime="10:38" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40324" daytime="10:39" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40325" daytime="10:40" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40326" daytime="10:41" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40327" daytime="10:42" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40328" daytime="10:43" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40329" daytime="10:44" number="18" order="18" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33693" />
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1297" daytime="10:45" gender="M" number="26" order="4" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1298" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1299" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1300" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1301" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1302" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1303" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1304" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1305" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1306" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40331" daytime="10:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40332" daytime="10:46" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40333" daytime="10:48" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40334" daytime="10:49" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40335" daytime="10:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40336" daytime="10:51" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40337" daytime="10:52" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40338" daytime="10:53" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40339" daytime="10:54" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40340" daytime="10:55" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40341" daytime="10:56" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40342" daytime="10:57" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40343" daytime="10:58" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40344" daytime="10:59" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40345" daytime="11:00" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40346" daytime="11:01" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40347" daytime="11:02" number="17" order="17" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1307" daytime="11:03" gender="F" number="27" order="5" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1308" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1309" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1310" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1311" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1312" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1313" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1314" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1315" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1316" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40348" daytime="11:03" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40349" daytime="11:07" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40350" daytime="11:11" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40351" daytime="11:15" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40352" daytime="11:18" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40353" daytime="11:22" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40354" daytime="11:25" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40355" daytime="11:29" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40356" daytime="11:32" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40357" daytime="11:35" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40358" daytime="11:39" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40359" daytime="11:42" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40360" daytime="11:45" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40361" daytime="11:48" number="14" order="14" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1317" daytime="11:51" gender="M" number="28" order="6" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1318" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1319" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1320" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1321" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1322" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1323" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1324" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1325" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1326" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40362" daytime="11:51" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40363" daytime="11:55" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40364" daytime="11:59" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40365" daytime="12:03" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40366" daytime="12:06" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40367" daytime="12:10" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40368" daytime="12:13" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40369" daytime="12:16" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40370" daytime="12:20" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40371" daytime="12:23" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40372" daytime="12:26" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40373" daytime="12:29" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40374" daytime="12:32" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40375" daytime="12:35" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40376" daytime="12:38" number="15" order="15" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1327" daytime="12:41" gender="F" number="29" order="7" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1328" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1329" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1330" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1331" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1332" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1333" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1334" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1335" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1336" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40377" daytime="12:41" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40378" daytime="12:44" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40379" daytime="12:46" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40380" daytime="12:48" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40381" daytime="12:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40382" daytime="12:52" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40383" daytime="12:54" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40384" daytime="12:56" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40385" daytime="12:58" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40386" daytime="13:00" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40387" daytime="13:02" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40388" daytime="13:04" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40389" daytime="13:06" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40390" daytime="13:08" number="14" order="14" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1337" daytime="13:10" gender="M" number="30" order="8" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1338" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1339" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1340" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1341" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1342" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1343" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1344" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1345" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1346" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40391" daytime="13:10" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40392" daytime="13:13" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40393" daytime="13:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40394" daytime="13:17" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40395" daytime="13:19" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40396" daytime="13:21" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40397" daytime="13:23" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40398" daytime="13:25" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40399" daytime="13:27" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40400" daytime="13:29" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40401" daytime="13:31" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40402" daytime="13:32" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40403" daytime="13:34" number="13" order="13" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2025-12-21" daytime="14:05" endtime="17:16" number="5" status="SEEDED">
          <EVENTS>
            <EVENT eventid="1347" daytime="14:05" gender="F" number="31" order="1" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1348" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1349" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1350" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1351" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1352" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1353" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1354" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1355" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1356" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40404" daytime="14:05" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40405" daytime="14:09" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40406" daytime="14:12" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40407" daytime="14:16" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40408" daytime="14:19" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40409" daytime="14:22" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40410" daytime="14:26" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40411" daytime="14:29" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40412" daytime="14:32" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40413" daytime="14:35" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40414" daytime="14:38" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40415" daytime="14:41" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40416" daytime="14:44" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40417" daytime="14:47" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40418" daytime="14:50" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40419" daytime="14:53" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40420" daytime="14:55" number="17" order="17" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1357" daytime="14:58" gender="M" number="32" order="2" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1358" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1359" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1360" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1361" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1362" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1363" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1364" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1365" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1366" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40421" daytime="14:58" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40422" daytime="15:02" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40423" daytime="15:06" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40424" daytime="15:09" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40425" daytime="15:12" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40426" daytime="15:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40427" daytime="15:18" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40428" daytime="15:22" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40429" daytime="15:25" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40430" daytime="15:27" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40431" daytime="15:30" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40432" daytime="15:33" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40433" daytime="15:36" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40434" daytime="15:39" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40435" daytime="15:41" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40436" daytime="15:44" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40437" daytime="15:47" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40438" daytime="15:49" number="18" order="18" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1367" daytime="15:52" gender="F" number="33" order="3" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1368" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1369" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1370" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1371" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1372" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1373" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1374" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1375" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1376" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40439" daytime="15:52" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40440" daytime="15:53" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40441" daytime="15:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40442" daytime="15:56" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40443" daytime="15:57" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40444" daytime="15:58" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40445" daytime="15:59" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40446" daytime="16:01" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40447" daytime="16:02" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40448" daytime="16:03" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40449" daytime="16:04" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40450" daytime="16:05" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40451" daytime="16:06" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40452" daytime="16:07" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40453" daytime="16:08" number="15" order="15" status="SEEDED" />
                <HEAT heatid="40454" daytime="16:10" number="16" order="16" status="SEEDED" />
                <HEAT heatid="40455" daytime="16:11" number="17" order="17" status="SEEDED" />
                <HEAT heatid="40456" daytime="16:12" number="18" order="18" status="SEEDED" />
                <HEAT heatid="40457" daytime="16:13" number="19" order="19" status="SEEDED" />
                <HEAT heatid="40458" daytime="16:14" number="20" order="20" status="SEEDED" />
                <HEAT heatid="40459" daytime="16:15" number="21" order="21" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1377" daytime="16:16" gender="M" number="34" order="4" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1378" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1379" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1380" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1381" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1382" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1383" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1384" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1385" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1386" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40460" daytime="16:16" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40461" daytime="16:18" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40462" daytime="16:19" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40463" daytime="16:20" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40464" daytime="16:21" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40465" daytime="16:22" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40466" daytime="16:23" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40467" daytime="16:25" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40468" daytime="16:26" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40469" daytime="16:27" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40470" daytime="16:28" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40471" daytime="16:29" number="12" order="12" status="SEEDED" />
                <HEAT heatid="40472" daytime="16:30" number="13" order="13" status="SEEDED" />
                <HEAT heatid="40473" daytime="16:31" number="14" order="14" status="SEEDED" />
                <HEAT heatid="40474" daytime="16:32" number="15" order="15" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1387" daytime="16:33" gender="F" number="35" order="5" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1388" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1389" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1390" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1391" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1392" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1393" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1394" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1395" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1396" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40475" daytime="16:33" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40476" daytime="16:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40477" daytime="16:38" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40478" daytime="16:40" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40479" daytime="16:42" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40480" daytime="16:43" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40481" daytime="16:45" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40482" daytime="16:47" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40483" daytime="16:49" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40484" daytime="16:51" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40485" daytime="16:52" number="11" order="11" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33677" />
                <TIMESTANDARDREF timestandardlistid="33679" />
                <TIMESTANDARDREF timestandardlistid="33681" />
                <TIMESTANDARDREF timestandardlistid="33683" />
                <TIMESTANDARDREF timestandardlistid="33685" />
                <TIMESTANDARDREF timestandardlistid="33687" />
                <TIMESTANDARDREF timestandardlistid="33689" />
                <TIMESTANDARDREF timestandardlistid="33691" />
                <TIMESTANDARDREF timestandardlistid="33693" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1397" daytime="16:54" gender="M" number="36" order="6" round="TIM" status="SEEDED" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE value="900" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1398" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1399" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1400" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1401" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1402" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1403" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1404" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1405" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1406" agemax="-1" agemin="18" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="40486" daytime="16:54" number="1" order="1" status="SEEDED" />
                <HEAT heatid="40487" daytime="16:56" number="2" order="2" status="SEEDED" />
                <HEAT heatid="40488" daytime="16:59" number="3" order="3" status="SEEDED" />
                <HEAT heatid="40489" daytime="17:01" number="4" order="4" status="SEEDED" />
                <HEAT heatid="40490" daytime="17:02" number="5" order="5" status="SEEDED" />
                <HEAT heatid="40491" daytime="17:04" number="6" order="6" status="SEEDED" />
                <HEAT heatid="40492" daytime="17:06" number="7" order="7" status="SEEDED" />
                <HEAT heatid="40493" daytime="17:08" number="8" order="8" status="SEEDED" />
                <HEAT heatid="40494" daytime="17:09" number="9" order="9" status="SEEDED" />
                <HEAT heatid="40495" daytime="17:11" number="10" order="10" status="SEEDED" />
                <HEAT heatid="40496" daytime="17:12" number="11" order="11" status="SEEDED" />
                <HEAT heatid="40497" daytime="17:14" number="12" order="12" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="33676" />
                <TIMESTANDARDREF timestandardlistid="33678" />
                <TIMESTANDARDREF timestandardlistid="33680" />
                <TIMESTANDARDREF timestandardlistid="33682" />
                <TIMESTANDARDREF timestandardlistid="33684" />
                <TIMESTANDARDREF timestandardlistid="33686" />
                <TIMESTANDARDREF timestandardlistid="33688" />
                <TIMESTANDARDREF timestandardlistid="33690" />
                <TIMESTANDARDREF timestandardlistid="33692" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="00883" nation="ESP" clubid="36951" name="Club Natación Calvià">
          <ATHLETES>
            <ATHLETE firstname="Adam " lastname="Tischer Rodríguez" birthdate="2013-01-01" gender="M" nation="ESP" license="1200426" athleteid="36952">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.33" eventid="1297" heatid="40333" lane="4" />
                <ENTRY entrytime="00:02:59.80" eventid="1317" heatid="40365" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5502" nation="GER" region="08" clubid="38862" name="Hanse SV Rostock">
          <ATHLETES>
            <ATHLETE firstname="Theodor" lastname="Rollow" birthdate="2005-01-01" gender="M" nation="GER" license="333696" athleteid="38863">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.35" eventid="1297" heatid="40345" lane="6">
                  <MEETINFO name="XIX. Rostock Masters Sprint Cup" city="Rostock" course="SCM" approved="GER" date="2025-06-21" qualificationtime="00:00:28.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.50" eventid="1377" heatid="40472" lane="3">
                  <MEETINFO name="XIX. Rostock Masters Sprint Cup" city="Rostock" course="SCM" approved="GER" date="2025-06-21" qualificationtime="00:00:29.84" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3358" nation="GER" region="12" clubid="38246" name="SWV TuR Dresden">
          <ATHLETES>
            <ATHLETE firstname="Lennox" lastname="Fischer" birthdate="2012-01-01" gender="M" nation="GER" license="445086" athleteid="38249">
              <ENTRIES>
                <ENTRY entrytime="00:09:46.84" eventid="1093" heatid="40017" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:09:46.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.40" eventid="1153" heatid="40109" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:37.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.52" eventid="1217" heatid="40185" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:34.66" />
                </ENTRY>
                <ENTRY entrytime="00:04:46.55" eventid="1257" heatid="40256" lane="1">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:04:46.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.07" eventid="1277" heatid="40299" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:02.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.40" eventid="1337" heatid="40400" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:13.80" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.75" eventid="1357" heatid="40432" lane="2">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:02:16.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Domke" birthdate="2009-01-01" gender="F" nation="GER" license="396910" athleteid="38247">
              <ENTRIES>
                <ENTRY entrytime="00:10:15.00" eventid="1083" heatid="40010" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Franka" lastname="Lukoschat" birthdate="2014-01-01" gender="F" nation="GER" license="458407" athleteid="38257">
              <ENTRIES>
                <ENTRY entrytime="00:11:30.60" eventid="1083" heatid="40005" lane="8" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4296" nation="GER" region="02" clubid="34621" name="SC Wfr. München">
          <ATHLETES>
            <ATHLETE firstname="Elias" lastname="Henkel" birthdate="2015-01-01" gender="M" nation="GER" license="461538" athleteid="37002">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.31" eventid="1133" heatid="40060" lane="6">
                  <MEETINFO name="49. Landshuter Pokalschwimmen" city="Landshut" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:38.04" />
                </ENTRY>
                <ENTRY entrytime="00:03:28.99" eventid="1173" heatid="40128" lane="7" />
                <ENTRY entrytime="00:00:46.40" eventid="1217" heatid="40175" lane="4">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:00:45.61" />
                </ENTRY>
                <ENTRY entrytime="00:06:12.99" eventid="1257" heatid="40246" lane="5">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:06:31.52" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.96" eventid="1297" heatid="40332" lane="7">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:41.96" />
                </ENTRY>
                <ENTRY entrytime="00:03:12.51" eventid="1317" heatid="40363" lane="5">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:03:09.37" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.63" eventid="1337" heatid="40393" lane="1">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:01:37.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Theodor" lastname="Engelmann" birthdate="2015-01-01" gender="M" nation="GER" license="464839" athleteid="36995">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.87" eventid="1133" heatid="40062" lane="7">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:35.33" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.62" eventid="1173" heatid="40131" lane="6">
                  <MEETINFO name="47. Internationales Feuerbacher Herbstschwimmen" city="Stuttgart" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:03:00.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.68" eventid="1237" heatid="40220" lane="1">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:01:21.29" />
                </ENTRY>
                <ENTRY entrytime="00:06:07.24" eventid="1257" heatid="40246" lane="4">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:06:07.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.46" eventid="1277" heatid="40291" lane="7">
                  <MEETINFO name="47. Internationales Feuerbacher Herbstschwimmen" city="Stuttgart" course="LCM" approved="GER" date="2025-11-16" qualificationtime="00:01:17.46" />
                </ENTRY>
                <ENTRY entrytime="00:03:20.62" eventid="1317" heatid="40362" lane="3">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:03:20.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Katharina" lastname="Schmidt" birthdate="2013-01-01" gender="F" nation="GER" license="497256" athleteid="37017">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.99" eventid="1267" heatid="40263" lane="4">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:18.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.99" eventid="1287" heatid="40313" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:00:39.69" />
                </ENTRY>
                <ENTRY entrytime="00:03:02.17" eventid="1347" heatid="40405" lane="7">
                  <MEETINFO name="28. Internationales Schwimmfest" city="München Obergiesing" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:58.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.96" eventid="1367" heatid="40441" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:41.96" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maximilian" lastname="Tack" birthdate="2014-01-01" gender="M" nation="GER" license="449444" athleteid="37032">
              <ENTRIES>
                <ENTRY entrytime="00:22:18.38" eventid="1113" heatid="40022" lane="6">
                  <MEETINFO name="Bay. Meisterschaften Lange Strecken" city="Würzburg" course="LCM" approved="GER" date="2025-01-18" qualificationtime="00:22:18.38" />
                </ENTRY>
                <ENTRY entrytime="00:03:15.48" eventid="1153" heatid="40104" lane="6">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:03:12.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.30" eventid="1173" heatid="40135" lane="7">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:02:47.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.67" eventid="1217" heatid="40178" lane="2">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:42.67" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.32" eventid="1237" heatid="40223" lane="1">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:01:19.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.53" eventid="1277" heatid="40293" lane="5">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:11.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.39" eventid="1337" heatid="40394" lane="3">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:28.87" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.98" eventid="1357" heatid="40424" lane="4">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:02:38.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.13" eventid="1377" heatid="40465" lane="7">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:37.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Johannes" lastname="Nibler" birthdate="2014-01-01" gender="M" nation="GER" license="451233" athleteid="37010">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.60" eventid="1133" heatid="40062" lane="2">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:35.60" />
                </ENTRY>
                <ENTRY entrytime="00:03:39.99" eventid="1197" heatid="40151" lane="3" />
                <ENTRY entrytime="00:05:58.65" eventid="1257" heatid="40247" lane="7">
                  <MEETINFO name="36. Int. Langstreckenschwimmen" city="Rosenheim" course="LCM" approved="GER" date="2025-06-01" qualificationtime="00:05:58.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.28" eventid="1277" heatid="40289" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:19.04" />
                </ENTRY>
                <ENTRY entrytime="00:03:17.24" eventid="1317" heatid="40362" lane="4">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:03:16.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.91" eventid="1357" heatid="40423" lane="6">
                  <MEETINFO name="36. Int. Langstreckenschwimmen" city="Rosenheim" course="LCM" approved="GER" date="2025-05-31" qualificationtime="00:02:50.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Quentin" lastname="Domurado" birthdate="2015-01-01" gender="M" nation="FRA" license="467535" athleteid="36986">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.18" eventid="1133" heatid="40060" lane="3">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:37.49" />
                </ENTRY>
                <ENTRY entrytime="00:03:40.99" eventid="1153" heatid="40102" lane="2">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:03:35.31" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.84" eventid="1237" heatid="40215" lane="3">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:32.89" />
                </ENTRY>
                <ENTRY entrytime="00:06:06.18" eventid="1257" heatid="40247" lane="8">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-18" qualificationtime="00:06:06.18" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.06" eventid="1277" heatid="40288" lane="4">
                  <MEETINFO name="36. Int. Langstreckenschwimmen" city="Rosenheim" course="LCM" approved="GER" date="2025-06-01" qualificationtime="00:01:21.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:47.68" eventid="1337" heatid="40391" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:46.72" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.06" eventid="1357" heatid="40422" lane="1">
                  <MEETINFO name="International Swim Meeting" city="Erlangen" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:02:59.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.16" eventid="1397" heatid="40487" lane="3">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:31.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Eva" lastname="Schreiner" birthdate="2012-01-01" gender="F" nation="GER" license="420331" athleteid="37022">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.87" eventid="1123" heatid="40041" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:31.87" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.94" eventid="1163" heatid="40117" lane="4">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:02:54.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.27" eventid="1227" heatid="40202" lane="2">
                  <MEETINFO name="28. Internationales Schwimmfest" city="München Obergiesing" course="SCM" approved="GER" date="2025-05-11" qualificationtime="00:01:17.56" />
                </ENTRY>
                <ENTRY entrytime="00:05:16.92" eventid="1247" heatid="40240" lane="7">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:05:16.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.43" eventid="1267" heatid="40276" lane="4">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:01:08.43" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.57" eventid="1307" heatid="40353" lane="8">
                  <MEETINFO name="47. Internationales Feuerbacher Herbstschwimmen" city="Stuttgart" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:02:49.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.38" eventid="1347" heatid="40415" lane="4">
                  <MEETINFO name="47. Internationales Feuerbacher Herbstschwimmen" city="Stuttgart" course="LCM" approved="GER" date="2025-11-16" qualificationtime="00:02:27.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paula" lastname="Seiwert" birthdate="2015-01-01" gender="F" nation="GER" license="470828" athleteid="37030" />
            <ATHLETE firstname="Theresa" lastname="Bär" birthdate="2015-01-01" gender="F" nation="GER" license="479601" athleteid="36978">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.50" eventid="1123" heatid="40027" lane="1">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:35.75" />
                </ENTRY>
                <ENTRY entrytime="00:03:32.32" eventid="1143" heatid="40091" lane="1">
                  <MEETINFO name="47. Internationales Feuerbacher Herbstschwimmen" city="Stuttgart" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:03:32.32" />
                </ENTRY>
                <ENTRY entrytime="00:06:13.99" eventid="1247" heatid="40234" lane="3" />
                <ENTRY entrytime="00:01:20.35" eventid="1267" heatid="40263" lane="3">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:01:17.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.41" eventid="1327" heatid="40379" lane="5">
                  <MEETINFO name="47. Internationales Feuerbacher Herbstschwimmen" city="Stuttgart" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:40.41" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.69" eventid="1347" heatid="40406" lane="3">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:02:48.71" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.99" eventid="1387" heatid="40476" lane="7" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Gabor" gender="M" lastname="Bordas" />
            <COACH firstname="Niklas" gender="M" lastname="Bressler" />
            <COACH firstname="Gabor" gender="M" lastname="Bordas" />
            <COACH firstname="Niklas" gender="M" lastname="Bressler" />
            <COACH firstname="Angela" gender="M" lastname="Leheis" />
            <COACH firstname="Angela" gender="M" lastname="Leheis" />
            <COACH firstname="Angela" gender="M" lastname="Leheis" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="4387" nation="GER" region="02" clubid="35622" name="SV Weiden">
          <ATHLETES>
            <ATHLETE firstname="Kira" lastname="Krawchina" birthdate="2013-01-01" gender="F" nation="GER" license="481523" athleteid="35677">
              <ENTRIES>
                <ENTRY entrytime="00:03:40.77" eventid="1143" heatid="40090" lane="2">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:03:40.77" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.99" eventid="1207" heatid="40159" lane="6">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:00:46.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.57" eventid="1267" heatid="40264" lane="2">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:19.42" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.00" eventid="1347" heatid="40405" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:03:02.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Friedrich" birthdate="2013-01-01" gender="M" nation="GER" license="445668" athleteid="35653">
              <ENTRIES>
                <ENTRY entrytime="00:02:58.90" eventid="1153" heatid="40107" lane="8">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:50.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.00" eventid="1217" heatid="40181" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:35.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.26" eventid="1297" heatid="40336" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:00:33.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.84" eventid="1337" heatid="40397" lane="3">
                  <MEETINFO name="8. Internationales Herbstmeeting" city="Mühlacker" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:18.38" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.00" eventid="1397" heatid="40488" lane="4">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:16.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leni" lastname="Dippold" birthdate="2009-01-01" gender="F" nation="GER" license="402050" athleteid="35641">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.65" eventid="1123" heatid="40051" lane="4">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:29.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.31" eventid="1267" heatid="40281" lane="4">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:03.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.52" eventid="1287" heatid="40327" lane="8">
                  <MEETINFO name="2. Int. Gugl Sprint Meeting" city="Linz" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:00:31.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.40" eventid="1387" heatid="40483" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:12.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Seidl" birthdate="2012-01-01" gender="M" nation="GER" license="441391" athleteid="35694">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.16" eventid="1133" heatid="40072" lane="3">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:29.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.86" eventid="1217" heatid="40179" lane="1">
                  <MEETINFO name="10. Kulmbacher Kinder-Schwimm-Vergnügen" city="Kulmbach" course="SCM" approved="GER" date="2025-02-22" qualificationtime="00:00:41.67" />
                </ENTRY>
                <ENTRY entrytime="00:05:10.00" eventid="1257" heatid="40253" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:05:00.77" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.02" eventid="1277" heatid="40298" lane="2">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:03.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.54" eventid="1337" heatid="40396" lane="1">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:25.60" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.70" eventid="1357" heatid="40428" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:20.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.88" eventid="1377" heatid="40464" lane="5">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:00:36.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Güll" birthdate="2006-01-01" gender="M" nation="GER" license="356936" athleteid="35665">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.98" eventid="1133" heatid="40086" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:25.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.37" eventid="1217" heatid="40186" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:00:34.15" />
                </ENTRY>
                <ENTRY entrytime="00:04:40.50" eventid="1257" heatid="40257" lane="6">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:04:44.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.54" eventid="1277" heatid="40310" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:00:55.81" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.80" eventid="1357" heatid="40436" lane="5">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:06.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nadja" lastname="Valea" birthdate="2007-01-01" gender="F" nation="GER" license="366678" athleteid="35718">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.04" eventid="1123" heatid="40057" lane="8">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:27.11" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.30" eventid="1267" heatid="40285" lane="3">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:00.11" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.54" eventid="1307" heatid="40358" lane="3">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:39.54" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jonas" lastname="Rupprecht" birthdate="2008-01-01" gender="M" nation="GER" license="425435" athleteid="35682">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.08" eventid="1133" heatid="40082" lane="6">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:26.66" />
                </ENTRY>
                <ENTRY entrytime="00:04:40.00" eventid="1257" heatid="40257" lane="5" />
                <ENTRY entrytime="00:01:00.42" eventid="1277" heatid="40305" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:57.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.62" eventid="1297" heatid="40342" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:29.44" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.00" eventid="1357" heatid="40432" lane="3">
                  <MEETINFO name="8. Internationales Herbstmeeting" city="Mühlacker" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:02:10.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Charlotte" lastname="Güll" birthdate="2009-01-01" gender="F" nation="GER" license="396729" athleteid="35659">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.54" eventid="1123" heatid="40055" lane="4">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:28.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.57" eventid="1207" heatid="40173" lane="7">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:34.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.55" eventid="1267" heatid="40284" lane="2">
                  <MEETINFO name="8. Internationales Herbstmeeting" city="Mühlacker" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:01.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.59" eventid="1287" heatid="40324" lane="3">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:00:32.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.45" eventid="1327" heatid="40390" lane="1">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:18.09" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Staeck" birthdate="2009-01-01" gender="F" nation="GER" license="497669" athleteid="35702">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.99" eventid="1123" heatid="40040" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:32.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.99" eventid="1227" heatid="40202" lane="6">
                  <MEETINFO name="10. Kulmbacher Kinder-Schwimm-Vergnügen" city="Kulmbach" course="SCM" approved="GER" date="2025-02-22" qualificationtime="00:01:21.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.50" eventid="1287" heatid="40319" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:35.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.62" eventid="1367" heatid="40449" lane="4">
                  <MEETINFO name="8. Internationales Herbstmeeting" city="Mühlacker" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:36.72" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Bauer" birthdate="2015-01-01" gender="F" nation="GER" license="471959" athleteid="35629">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.09" eventid="1123" heatid="40029" lane="4">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:00:34.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.69" eventid="1227" heatid="40195" lane="2">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:29.17" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.71" eventid="1267" heatid="40264" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:15.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.39" eventid="1287" heatid="40312" lane="1">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:00:37.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.55" eventid="1367" heatid="40443" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:38.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anton" lastname="Seidl" birthdate="2014-01-01" gender="M" nation="GER" license="454046" athleteid="35688">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.33" eventid="1133" heatid="40060" lane="2">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:36.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.83" eventid="1217" heatid="40175" lane="6">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:46.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.64" eventid="1277" heatid="40289" lane="1">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:20.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:42.34" eventid="1337" heatid="40392" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:42.34" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.77" eventid="1357" heatid="40422" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:03:02.07" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Frida" lastname="Wegerer" birthdate="2011-01-01" gender="F" nation="GER" license="479924" athleteid="35722">
              <ENTRIES>
                <ENTRY entrytime="00:11:00.00" eventid="1083" heatid="40007" lane="3" />
                <ENTRY entrytime="00:00:31.90" eventid="1123" heatid="40040" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:30.56" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.06" eventid="1247" heatid="40240" lane="5">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:05:15.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.81" eventid="1267" heatid="40275" lane="4">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:06.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.50" eventid="1327" heatid="40382" lane="3">
                  <MEETINFO name="10. Kulmbacher Kinder-Schwimm-Vergnügen" city="Kulmbach" course="SCM" approved="GER" date="2025-02-22" qualificationtime="00:01:32.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.00" eventid="1347" heatid="40411" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:27.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Friedrich" birthdate="2014-01-01" gender="F" nation="GER" license="454047" athleteid="35646">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.00" eventid="1123" heatid="40026" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:37.96" />
                </ENTRY>
                <ENTRY entrytime="00:03:45.00" eventid="1143" heatid="40090" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:03:50.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.50" eventid="1207" heatid="40158" lane="1">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:49.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.53" eventid="1267" heatid="40262" lane="2">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:23.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.99" eventid="1327" heatid="40378" lane="6">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:48.17" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.00" eventid="1347" heatid="40406" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:56.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Andrey" lastname="Klein" birthdate="2014-01-01" gender="M" nation="GER" license="481516" athleteid="35671">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.42" eventid="1133" heatid="40062" lane="3">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:00:33.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.81" eventid="1217" heatid="40176" lane="7">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:00:45.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.98" eventid="1277" heatid="40289" lane="8">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:15.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.48" eventid="1337" heatid="40392" lane="5">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:39.61" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.00" eventid="1357" heatid="40422" lane="5">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:49.23" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Victoria-Sophia" lastname="Titz" birthdate="2015-01-01" gender="F" nation="GER" license="471957" athleteid="35712">
              <ENTRIES>
                <ENTRY entrytime="00:03:16.09" eventid="1163" heatid="40113" lane="6">
                  <MEETINFO name="12. BSV Bezirksvergleich im Schwimmen" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:03:13.91" />
                </ENTRY>
                <ENTRY entrytime="00:06:15.99" eventid="1247" heatid="40233" lane="4">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:06:35.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.00" eventid="1267" heatid="40261" lane="5">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:01:26.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.81" eventid="1327" heatid="40378" lane="1">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:45.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.70" eventid="1367" heatid="40440" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:43.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sina" lastname="Strohmeier" birthdate="2010-01-01" gender="F" nation="GER" license="457642" athleteid="35707">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.18" eventid="1123" heatid="40035" lane="1">
                  <MEETINFO name="8. Internationales Herbstmeeting" city="Mühlacker" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:33.21" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.99" eventid="1267" heatid="40271" lane="4">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:14.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.50" eventid="1287" heatid="40315" lane="6">
                  <MEETINFO name="24. Kurfürstenpokal Amberg" city="Amberg" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:00:37.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.50" eventid="1367" heatid="40446" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:40.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hannah" lastname="Bauer" birthdate="2012-01-01" gender="F" nation="GER" license="454444" athleteid="35623">
              <ENTRIES>
                <ENTRY entrytime="00:05:50.99" eventid="1063" heatid="39995" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:06:12.34" />
                </ENTRY>
                <ENTRY entrytime="00:03:25.00" eventid="1143" heatid="40092" lane="1">
                  <MEETINFO name="8. Internationales Herbstmeeting" city="Mühlacker" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:03:19.78" />
                </ENTRY>
                <ENTRY entrytime="00:03:15.00" eventid="1187" heatid="40147" lane="3">
                  <MEETINFO name="8. Internationales Herbstmeeting" city="Mühlacker" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:03:09.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.20" eventid="1287" heatid="40314" lane="6">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:37.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.00" eventid="1387" heatid="40478" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:21.49" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emma" lastname="Wutz" birthdate="2008-01-01" gender="F" nation="GER" license="370566" athleteid="35729">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.03" eventid="1123" heatid="40045" lane="5">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:30.38" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.07" eventid="1267" heatid="40275" lane="5">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:07.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.00" eventid="1287" heatid="40318" lane="1">
                  <MEETINFO name="2. Int. Gugl Sprint Meeting" city="Linz" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:00:35.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.19" eventid="1367" heatid="40448" lane="5">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:37.19" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marie" lastname="Binner" birthdate="2012-01-01" gender="F" nation="GER" license="441395" athleteid="35635">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.74" eventid="1123" heatid="40036" lane="2">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:00:32.74" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.83" eventid="1163" heatid="40116" lane="1">
                  <MEETINFO name="DMS-Austragung 24/25 Bezirksliga - Oberpfalz" city="Weiden" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:02:58.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.29" eventid="1227" heatid="40199" lane="3">
                  <MEETINFO name="30. Internationales Adventspokalschwimmen" city="Tirschenreuth" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:21.33" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.00" eventid="1307" heatid="40350" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:02:58.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.00" eventid="1367" heatid="40447" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:37.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:16.00" eventid="1185" heatid="40145" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="35682" number="1" />
                    <RELAYPOSITION athleteid="35653" number="2" />
                    <RELAYPOSITION athleteid="35694" number="3" />
                    <RELAYPOSITION athleteid="35665" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" date="2025-11-15" qualificationtime="00:02:16.50" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:17.00" eventid="1183" heatid="40143" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="35729" number="1" />
                    <RELAYPOSITION athleteid="35718" number="2" />
                    <RELAYPOSITION athleteid="35641" number="3" />
                    <RELAYPOSITION athleteid="35707" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="8. Internationales Herbstmeeting" city="Mühlacker" date="2025-11-02" qualificationtime="00:02:20.51" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4292" nation="GER" region="02" clubid="34858" name="SC Prinz Eugen München">
          <ATHLETES>
            <ATHLETE firstname="Lea" lastname="Czeczko" birthdate="2008-01-01" gender="F" nation="GER" license="377570" athleteid="34859">
              <ENTRIES>
                <ENTRY entrytime="00:05:47.34" eventid="1063" heatid="39996" lane="1">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:05:47.34" />
                </ENTRY>
                <ENTRY entrytime="00:11:00.59" eventid="1083" heatid="40007" lane="6" />
                <ENTRY entrytime="00:03:08.52" eventid="1143" heatid="40095" lane="1" />
                <ENTRY entrytime="00:02:43.04" eventid="1163" heatid="40122" lane="4">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-10" qualificationtime="00:02:43.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.41" eventid="1207" heatid="40162" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Mangafic" gender="M" lastname="Elvir - Elli" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" clubid="34688" name="Kampfrichter">
          <OFFICIALS>
            <OFFICIAL officialid="52" firstname="Maja" gender="F" lastname="Neubert" />
            <OFFICIAL officialid="39" firstname="Paul" gender="M" lastname="Leinung" />
            <OFFICIAL officialid="22" firstname="Nathalie" gender="F" lastname="Grohneberg" />
            <OFFICIAL officialid="1" firstname="Antje" gender="F" lastname="Abraham" />
            <OFFICIAL officialid="82" firstname="Andreas" gender="M" lastname="Trodler" />
            <OFFICIAL officialid="77" firstname="Matthias" gender="M" lastname="Schubert" />
            <OFFICIAL officialid="14643" firstname="Niclas" gender="M" lastname="Lang" />
            <OFFICIAL officialid="20601" firstname="Oliver" gender="M" lastname="Otti" />
            <OFFICIAL officialid="55" firstname="Falk" gender="M" lastname="Nietsch" />
            <OFFICIAL officialid="38" firstname="Martina" gender="F" lastname="Lehnhardt" />
            <OFFICIAL officialid="17" firstname="Ricarda" gender="F" lastname="Forkert" />
            <OFFICIAL officialid="98" firstname="Markus" gender="M" lastname="Zomack" />
            <OFFICIAL officialid="93" firstname="Tom" gender="M" lastname="Wiedemann" />
            <OFFICIAL officialid="76" firstname="Cornelius" gender="M" lastname="Schramm" />
            <OFFICIAL officialid="20602" firstname="Julian Alexander" gender="M" lastname="Nietzold" />
            <OFFICIAL officialid="5998" firstname="Anika" gender="F" lastname="Böhme" />
            <OFFICIAL officialid="54" firstname="Sina" gender="F" lastname="Neumeister" />
            <OFFICIAL officialid="33" firstname="Franziska" gender="F" lastname="Kionke" />
            <OFFICIAL officialid="16" firstname="Robin" gender="M" lastname="Erdmann" />
            <OFFICIAL officialid="3" firstname="Gregor" gender="M" lastname="Abraham" />
            <OFFICIAL officialid="92" firstname="Ute" gender="F" lastname="Weinhold" />
            <OFFICIAL officialid="79" firstname="Olaf" gender="M" lastname="Schulz" />
            <OFFICIAL officialid="36007" firstname="Birgit" gender="F" lastname="Beckmann" />
            <OFFICIAL officialid="20596" firstname="Doreen" gender="F" lastname="Barthel" />
            <OFFICIAL officialid="49" firstname="Marie" gender="F" lastname="Müller" />
            <OFFICIAL officialid="32" firstname="Gesa Luise" gender="F" lastname="Kempe" />
            <OFFICIAL officialid="19" firstname="Fabian" gender="M" lastname="Gärtner" />
            <OFFICIAL officialid="2" firstname="Peter" gender="M" lastname="Abraham" />
            <OFFICIAL officialid="5949" firstname="Pauline" gender="F" lastname="Markert" />
            <OFFICIAL officialid="5937" firstname="Sophia" gender="F" lastname="Lorenz" />
            <OFFICIAL officialid="95" firstname="Tom" gender="M" lastname="Wiese" />
            <OFFICIAL officialid="78" firstname="Reinhard" gender="M" lastname="Schultz" />
            <OFFICIAL officialid="14606" firstname="Alexander" gender="M" lastname="Beier" />
            <OFFICIAL officialid="20594" firstname="Lars" gender="M" lastname="Martin" />
            <OFFICIAL officialid="35859" firstname="Maren" gender="F" lastname="Böhme" />
            <OFFICIAL officialid="14585" firstname="Uwe" gender="M" lastname="Albert" />
            <OFFICIAL officialid="48" firstname="Anton" gender="M" lastname="Müller" />
            <OFFICIAL officialid="35" firstname="Maria" gender="F" lastname="Küllig" />
            <OFFICIAL officialid="18" firstname="Thomas" gender="M" lastname="Funke" />
            <OFFICIAL officialid="13" firstname="Sandra" gender="F" lastname="Conseur" />
            <OFFICIAL officialid="14610" firstname="Liam" gender="M" lastname="Rühmann" />
            <OFFICIAL officialid="35865" firstname="Steffen" gender="M" lastname="Böhmert" />
            <OFFICIAL officialid="94" firstname="Manja" gender="F" lastname="Wiese" />
            <OFFICIAL officialid="73" firstname="Tim" gender="M" lastname="Schneider" />
            <OFFICIAL officialid="5930" firstname="Jens" gender="M" lastname="Böhmert" />
            <OFFICIAL officialid="14594" firstname="Nadine" gender="F" lastname="Engmann" />
            <OFFICIAL officialid="51" firstname="Eileen" gender="F" lastname="Neubert" />
            <OFFICIAL officialid="34" firstname="Christina" gender="F" lastname="Knorr" />
            <OFFICIAL officialid="29" firstname="Ina" gender="F" lastname="Humburg" />
            <OFFICIAL officialid="12" firstname="Jan" gender="M" lastname="Böhmert" />
            <OFFICIAL officialid="20604" firstname="Manuela" gender="F" lastname="Seibel" />
            <OFFICIAL officialid="20606" firstname="Martin" gender="M" lastname="Kupfer" />
            <OFFICIAL officialid="89" firstname="Rika" gender="F" lastname="Wappler" />
            <OFFICIAL officialid="72" firstname="Frank" gender="M" lastname="Schmiedel" />
            <OFFICIAL officialid="35862" firstname="Leonie" gender="F" lastname="Wiese" />
            <OFFICIAL officialid="35864" firstname="Lilo" gender="F" lastname="Firkert" />
            <OFFICIAL officialid="14683" firstname="Judith" gender="F" lastname="Schreiber" />
            <OFFICIAL officialid="5935" firstname="Sabine" gender="F" lastname="Eder" />
            <OFFICIAL officialid="36005" firstname="Thomwas" gender="M" lastname="Werdin" />
            <OFFICIAL officialid="50" firstname="Susann" gender="F" lastname="Naumann" />
            <OFFICIAL officialid="45" firstname="Sonja" gender="F" lastname="Mehnert" />
            <OFFICIAL officialid="28" firstname="Malte" gender="M" lastname="Hoffbauer" />
            <OFFICIAL officialid="15" firstname="Maximilian" gender="M" lastname="Eichelkraut" />
            <OFFICIAL officialid="88" firstname="Mirko" gender="M" lastname="Wappler" />
            <OFFICIAL officialid="75" firstname="Sandro" gender="M" lastname="Schoop" />
            <OFFICIAL officialid="5944" firstname="Theresa" gender="F" lastname="Freytag" />
            <OFFICIAL officialid="36004" firstname="Severine" gender="F" lastname="Banek" />
            <OFFICIAL officialid="61" firstname="Sarah" gender="F" lastname="Rößler" />
            <OFFICIAL officialid="44" firstname="Thomas" gender="M" lastname="Medack" />
            <OFFICIAL officialid="31" firstname="Birgit" gender="F" lastname="Kaiser" />
            <OFFICIAL officialid="14" firstname="Alexa" gender="F" lastname="Ehrentraut" />
            <OFFICIAL officialid="91" firstname="Steffen" gender="M" lastname="Wegner" />
            <OFFICIAL officialid="74" firstname="Jeannette" gender="F" lastname="Schönherr" />
            <OFFICIAL officialid="69" firstname="André" gender="M" lastname="Schlott" />
            <OFFICIAL officialid="36002" firstname="Pepe" gender="M" lastname="Tzschoppe" />
            <OFFICIAL officialid="20595" firstname="Jens" gender="M" lastname="Fähndrich" />
            <OFFICIAL officialid="60" firstname="Lara Marie" gender="F" lastname="Peter" />
            <OFFICIAL officialid="47" firstname="Alexander" gender="M" lastname="Müller" />
            <OFFICIAL officialid="30" firstname="Hannah" gender="F" lastname="Johne" />
            <OFFICIAL officialid="9" firstname="Katrin" gender="F" lastname="Bodusch" />
            <OFFICIAL officialid="20712" firstname="Niclas" gender="M" lastname="Kühn" />
            <OFFICIAL officialid="90" firstname="Carina" gender="F" lastname="Wegner" />
            <OFFICIAL officialid="85" firstname="Jörg" gender="M" lastname="Volejnik" />
            <OFFICIAL officialid="68" firstname="Matthias" gender="M" lastname="Schliesch" />
            <OFFICIAL officialid="14590" firstname="Roy" gender="M" lastname="Wachsmuth" />
            <OFFICIAL officialid="20668" firstname="Martin" gender="M" lastname="Jähnel" />
            <OFFICIAL officialid="63" firstname="André" gender="M" lastname="Sauer" />
            <OFFICIAL officialid="46" firstname="Claudia" gender="F" lastname="Menke" />
            <OFFICIAL officialid="25" firstname="Alix" gender="F" lastname="Günther" />
            <OFFICIAL officialid="8" firstname="Lars" gender="M" lastname="Bludau" />
            <OFFICIAL officialid="20670" firstname="Matthias" gender="M" lastname="Malecki" />
            <OFFICIAL officialid="35863" firstname="Andrea" gender="F" lastname="Kirberger " />
            <OFFICIAL officialid="36001" firstname="Daniel" gender="M" lastname="Bingenheimer" />
            <OFFICIAL officialid="71" firstname="Carolyn Christin" gender="F" lastname="Schmidt" />
            <OFFICIAL officialid="62" firstname="Silke" gender="F" lastname="Rößler" />
            <OFFICIAL officialid="41" firstname="Joshua" gender="M" lastname="Liebelt" />
            <OFFICIAL officialid="24" firstname="Thomas" gender="M" lastname="Große" />
            <OFFICIAL officialid="11" firstname="Sven" gender="M" lastname="Böhme" />
            <OFFICIAL officialid="14681" firstname="Emily" gender="M" lastname="Schulz" />
            <OFFICIAL officialid="20603" firstname="Stefanie" gender="F" lastname="Bethge" />
            <OFFICIAL officialid="14603" firstname="Jasmin" gender="F" lastname="Zesewitz" />
            <OFFICIAL officialid="87" firstname="Petra" gender="F" lastname="Volejnik" />
            <OFFICIAL officialid="70" firstname="Laura" gender="F" lastname="Schlott" />
            <OFFICIAL officialid="20711" firstname="Julia" gender="F" lastname="Jentzsch" />
            <OFFICIAL officialid="36000" firstname="Alexander" gender="M" lastname="Kral" />
            <OFFICIAL officialid="57" firstname="Antje" gender="F" lastname="Oehme" />
            <OFFICIAL officialid="40" firstname="Simon" gender="M" lastname="Lerche" />
            <OFFICIAL officialid="27" firstname="Benedict" gender="M" lastname="Hildesheim" />
            <OFFICIAL officialid="10" firstname="Elke" gender="F" lastname="Böhm" />
            <OFFICIAL officialid="5" firstname="Ines" gender="F" lastname="Beck" />
            <OFFICIAL officialid="5946" firstname="Julia" gender="F" lastname="Knott" />
            <OFFICIAL officialid="20597" firstname="Stephanie" gender="F" lastname="Schmidt" />
            <OFFICIAL officialid="86" firstname="Kai" gender="M" lastname="Volejnik" />
            <OFFICIAL officialid="65" firstname="Mandy" gender="F" lastname="Scheffler" />
            <OFFICIAL officialid="5933" firstname="Anett" gender="F" lastname="Jacob" />
            <OFFICIAL officialid="5954" firstname="Gabriela" gender="F" lastname="Harnisch" />
            <OFFICIAL officialid="20651" firstname="Ana" gender="F" lastname="Pasquali de Hallier" />
            <OFFICIAL officialid="14680" firstname="Kathleen" gender="F" lastname="Woßeng" />
            <OFFICIAL officialid="35866" firstname="Maika" gender="F" lastname="Przisambor" />
            <OFFICIAL officialid="36003" firstname="Pauline" gender="F" lastname="Kohl" />
            <OFFICIAL officialid="56" firstname="Uta" gender="F" lastname="Oehlert" />
            <OFFICIAL officialid="43" firstname="Beatrix" gender="F" lastname="Mahn" />
            <OFFICIAL officialid="26" firstname="Ulrich" gender="M" lastname="Henning" />
            <OFFICIAL officialid="21" firstname="Richard" gender="M" lastname="Grohmann" />
            <OFFICIAL officialid="4" firstname="Mick" gender="M" lastname="Balzer" />
            <OFFICIAL officialid="5993" firstname="Torsten" gender="M" lastname="Naumann" />
            <OFFICIAL officialid="20598" firstname="Antje" gender="F" lastname="Deichmüller" />
            <OFFICIAL officialid="81" firstname="Annika" gender="F" lastname="Stange" />
            <OFFICIAL officialid="64" firstname="Anne" gender="F" lastname="Sauer" />
            <OFFICIAL officialid="35861" firstname="Steffi" gender="F" lastname="Böhmert" />
            <OFFICIAL officialid="5959" firstname="Claus" gender="M" lastname="Franke" />
            <OFFICIAL officialid="59" firstname="Robin" gender="M" lastname="Oehme" />
            <OFFICIAL officialid="42" firstname="Sandra" gender="F" lastname="Liebs" />
            <OFFICIAL officialid="37" firstname="Andrea" gender="F" lastname="Langner" />
            <OFFICIAL officialid="20" firstname="Robin" gender="M" lastname="Goldberg" />
            <OFFICIAL officialid="7" firstname="Silvia" gender="F" lastname="Beutin" />
            <OFFICIAL officialid="20599" firstname="André" gender="M" lastname="Matthes" />
            <OFFICIAL officialid="97" firstname="Daniela" gender="F" lastname="Zische" />
            <OFFICIAL officialid="80" firstname="Oskar" gender="M" lastname="Schwamberger" />
            <OFFICIAL officialid="67" firstname="Svenja" gender="F" lastname="Schlicke" />
            <OFFICIAL officialid="5939" firstname="Oliver" gender="M" lastname="Haberkorn" />
            <OFFICIAL officialid="20672" firstname="Marie" gender="F" lastname="Kiefer" />
            <OFFICIAL officialid="35860" firstname="Caroline" gender="F" lastname="Schulze" />
            <OFFICIAL officialid="36006" firstname="Martin" gender="M" lastname="Sykora" />
            <OFFICIAL officialid="58" firstname="Dirk" gender="M" lastname="Oehme" />
            <OFFICIAL officialid="53" firstname="Susann" gender="F" lastname="Neumann" />
            <OFFICIAL officialid="36" firstname="Katrin" gender="F" lastname="Lange" />
            <OFFICIAL officialid="23" firstname="Carolin" gender="F" lastname="Groneberg" />
            <OFFICIAL officialid="6" firstname="Yvonne" gender="F" lastname="Beier" />
            <OFFICIAL officialid="35858" firstname="Sophia" gender="F" lastname="Beier" />
            <OFFICIAL officialid="96" firstname="Philipp" gender="M" lastname="Wollmann" />
            <OFFICIAL officialid="83" firstname="Marcus" gender="M" lastname="Ulbricht" />
            <OFFICIAL officialid="66" firstname="Michael" gender="M" lastname="Schellhammer" />
            <OFFICIAL officialid="35999" firstname="Louis Matthias" gender="M" lastname="Dietrich" />
            <OFFICIAL officialid="20600" firstname="Sophia" gender="F" lastname="Uschakow" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="ESAHK" nation="CZE" clubid="38984" name="Elite Standart Academy">
          <CONTACT country="CZ" name="Marek Kovar" />
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Kertész" birthdate="2009-01-01" gender="M" nation="CZE" athleteid="39007">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.90" eventid="1133" heatid="40080" lane="8">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:28.01" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.00" eventid="1153" heatid="40108" lane="1">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:52.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.00" eventid="1217" heatid="40185" lane="4">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:35.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.99" eventid="1277" heatid="40306" lane="7" />
                <ENTRY entrytime="00:00:29.00" eventid="1297" heatid="40343" lane="2">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:29.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.00" eventid="1337" heatid="40399" lane="4" />
                <ENTRY entrytime="00:02:12.00" eventid="1357" heatid="40434" lane="5">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:12.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.00" eventid="1377" heatid="40473" lane="3">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:31.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Vnuková" birthdate="2009-01-01" gender="F" nation="CZE" athleteid="39066">
              <ENTRIES>
                <ENTRY entrytime="00:10:00.00" eventid="1083" status="WDR" />
                <ENTRY entrytime="00:02:55.00" eventid="1143" status="WDR" />
                <ENTRY entrytime="00:00:39.00" eventid="1207" status="WDR" />
                <ENTRY entrytime="00:05:00.00" eventid="1247" status="WDR" />
                <ENTRY entrytime="00:01:04.00" eventid="1267" status="WDR">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:06.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.00" eventid="1307" status="WDR" />
                <ENTRY entrytime="00:02:20.00" eventid="1347" status="WDR">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:19.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.00" eventid="1387" status="WDR">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:12.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Kertész" birthdate="2012-01-01" gender="F" nation="CZE" athleteid="39026">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.00" eventid="1123" heatid="40050" lane="2">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:30.34" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.00" eventid="1143" heatid="40097" lane="5" />
                <ENTRY entrytime="00:03:15.00" eventid="1187" heatid="40147" lane="5" />
                <ENTRY entrytime="00:00:36.00" eventid="1207" heatid="40172" lane="5">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:36.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.00" eventid="1287" heatid="40323" lane="2">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.54" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.00" eventid="1307" heatid="40358" lane="2" />
                <ENTRY entrytime="00:02:20.00" eventid="1347" heatid="40418" lane="2" />
                <ENTRY entrytime="00:01:20.00" eventid="1387" heatid="40479" lane="7" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Matěj" lastname="Šmíd" birthdate="2012-01-01" gender="M" nation="CZE" athleteid="38995">
              <ENTRIES>
                <ENTRY entrytime="00:05:20.00" eventid="1073" heatid="40000" lane="4" />
                <ENTRY entrytime="00:09:36.00" eventid="1093" heatid="40017" lane="4" />
                <ENTRY entrytime="00:02:46.00" eventid="1153" heatid="40109" lane="7" />
                <ENTRY entrytime="00:02:32.00" eventid="1173" heatid="40138" lane="5" />
                <ENTRY entrytime="00:02:45.00" eventid="1197" heatid="40153" lane="3" />
                <ENTRY entrytime="00:04:44.00" eventid="1257" heatid="40256" lane="5" />
                <ENTRY entrytime="00:01:03.00" eventid="1277" heatid="40302" lane="2" />
                <ENTRY entrytime="00:00:31.00" eventid="1297" heatid="40340" lane="6" />
                <ENTRY entrytime="00:01:22.00" eventid="1337" heatid="40397" lane="5" />
                <ENTRY entrytime="00:02:13.00" eventid="1357" heatid="40434" lane="7" />
                <ENTRY entrytime="00:00:32.50" eventid="1377" heatid="40470" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karolína" lastname="Serbousková" birthdate="2012-01-01" gender="F" nation="CZE" athleteid="39035">
              <ENTRIES>
                <ENTRY entrytime="00:10:54.00" eventid="1083" heatid="40008" lane="1" />
                <ENTRY entrytime="00:00:32.00" eventid="1123" heatid="40039" lane="6">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:33.35" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.00" eventid="1163" heatid="40122" lane="2">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:44.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.00" eventid="1187" heatid="40149" lane="8">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:52.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.00" eventid="1227" heatid="40207" lane="2">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:16.71" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.00" eventid="1267" heatid="40277" lane="3">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:08.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.00" eventid="1287" heatid="40323" lane="7">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:35.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.00" eventid="1367" heatid="40451" lane="7">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:36.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.00" eventid="1387" heatid="40481" lane="6">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:19.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Veronika" lastname="Krejčíková" birthdate="2012-01-01" gender="F" nation="CZE" athleteid="39056">
              <ENTRIES>
                <ENTRY entrytime="00:11:45.00" eventid="1083" heatid="40004" lane="2" />
                <ENTRY entrytime="00:00:31.99" eventid="1123" heatid="40039" lane="5" />
                <ENTRY entrytime="00:02:58.00" eventid="1163" heatid="40116" lane="5" />
                <ENTRY entrytime="00:00:42.00" eventid="1207" heatid="40163" lane="8" />
                <ENTRY entrytime="00:01:23.00" eventid="1227" heatid="40200" lane="8">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:23.39" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.00" eventid="1267" heatid="40273" lane="7">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:10.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.00" eventid="1307" heatid="40352" lane="3">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:58.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.00" eventid="1347" heatid="40409" lane="5">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:41.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.99" eventid="1367" heatid="40447" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Zajíc" birthdate="2010-01-01" gender="M" nation="CZE" athleteid="39016">
              <ENTRIES>
                <ENTRY entrytime="00:05:20.00" eventid="1073" heatid="40001" lane="8" />
                <ENTRY entrytime="00:00:27.00" eventid="1133" heatid="40083" lane="2">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:27.19" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.00" eventid="1153" heatid="40109" lane="2" />
                <ENTRY entrytime="00:02:35.00" eventid="1197" heatid="40154" lane="2">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:31.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.99" eventid="1217" heatid="40187" lane="6">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:33.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.00" eventid="1297" heatid="40344" lane="5">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:28.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.00" eventid="1337" heatid="40401" lane="2" />
                <ENTRY entrytime="00:02:15.00" eventid="1357" heatid="40433" lane="8">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:13.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.00" eventid="1397" heatid="40494" lane="6">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:05.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Adéla" lastname="Novotná" birthdate="2013-01-01" gender="F" nation="CZE" athleteid="39045">
              <ENTRIES>
                <ENTRY entrytime="00:05:50.00" eventid="1063" heatid="39996" lane="8" />
                <ENTRY entrytime="00:00:30.00" eventid="1123" heatid="40050" lane="7">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:31.56" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.00" eventid="1143" heatid="40097" lane="8" />
                <ENTRY entrytime="00:00:40.00" eventid="1207" heatid="40166" lane="6">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:40.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.00" eventid="1227" heatid="40208" lane="6">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:15.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.00" eventid="1267" heatid="40281" lane="7">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:05.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.00" eventid="1287" heatid="40321" lane="8">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.80" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.00" eventid="1307" heatid="40357" lane="7">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:45.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.00" eventid="1367" heatid="40455" lane="3">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:36.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.00" eventid="1387" heatid="40480" lane="6">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:18.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Štěpán" lastname="Šmíd" birthdate="2014-01-01" gender="M" nation="CZE" athleteid="38985">
              <ENTRIES>
                <ENTRY entrytime="00:20:45.00" eventid="1113" heatid="40024" lane="8" />
                <ENTRY entrytime="00:00:31.00" eventid="1133" heatid="40071" lane="8" />
                <ENTRY entrytime="00:02:42.00" eventid="1173" heatid="40136" lane="2" />
                <ENTRY entrytime="00:00:40.00" eventid="1217" heatid="40179" lane="5" />
                <ENTRY entrytime="00:05:20.00" eventid="1257" heatid="40251" lane="3" />
                <ENTRY entrytime="00:00:33.00" eventid="1297" heatid="40337" lane="2" />
                <ENTRY entrytime="00:01:26.00" eventid="1337" heatid="40396" lane="5" />
                <ENTRY entrytime="00:02:30.00" eventid="1357" heatid="40428" lane="8" />
                <ENTRY entrytime="00:00:36.00" eventid="1377" heatid="40466" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6615" nation="GER" region="07" clubid="38176" name="VFS Rödermark">
          <ATHLETES>
            <ATHLETE firstname="Lisa" lastname="Schader" birthdate="2010-01-01" gender="F" nation="GER" license="409186" athleteid="38224">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.57" eventid="1123" heatid="40055" lane="5">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:28.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.74" eventid="1227" heatid="40212" lane="4">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:08.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.79" eventid="1287" heatid="40328" lane="5">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-23" qualificationtime="00:00:30.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.93" eventid="1367" heatid="40457" lane="3">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:32.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Schickedanz" birthdate="2011-01-01" gender="F" nation="GER" license="427170" athleteid="38229">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.63" eventid="1123" heatid="40033" lane="3">
                  <MEETINFO name="Bezirks- und Bezirksjahrgangsmeisterschaften" city="Darmstadt" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:00:33.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.66" eventid="1267" heatid="40265" lane="8">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:18.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.00" eventid="1287" heatid="40314" lane="3" />
                <ENTRY entrytime="00:00:42.80" eventid="1367" heatid="40440" lane="4">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:42.80" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Hofferbert" birthdate="2008-01-01" gender="F" nation="GER" license="387377" athleteid="38177">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.31" eventid="1123" heatid="40044" lane="3">
                  <MEETINFO name="BaHaMa Cup" city="Langen" course="LCM" approved="GER" date="2025-03-22" qualificationtime="00:00:31.31" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.98" eventid="1227" heatid="40203" lane="5">
                  <MEETINFO name="44. Drei-Länder-Pokal" city="Lampertheim" course="SCM" approved="GER" date="2025-03-09" qualificationtime="00:01:18.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.10" eventid="1267" heatid="40273" lane="8">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:09.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.63" eventid="1367" heatid="40448" lane="1">
                  <MEETINFO name="44. Drei-Länder-Pokal" city="Lampertheim" course="SCM" approved="GER" date="2025-03-09" qualificationtime="00:00:36.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Semih" lastname="Taskin" birthdate="2009-01-01" gender="M" nation="GER" license="399722" athleteid="38239">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.89" eventid="1133" heatid="40083" lane="5">
                  <MEETINFO name="Hochtaunus-Cup" city="Oberursel" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:26.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.69" eventid="1217" heatid="40187" lane="5">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:33.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.07" eventid="1277" heatid="40305" lane="5">
                  <MEETINFO name="Kreismeisterschaft Offenbach/Einlagungswettkampf" city="Heusenstamm" course="SCM" approved="GER" date="2025-11-29" qualificationtime="00:01:01.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.01" eventid="1337" heatid="40400" lane="1">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:14.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.46" eventid="1377" heatid="40469" lane="4">
                  <MEETINFO name="Kreismeisterschaft Offenbach/Einlagungswettkampf" city="Heusenstamm" course="SCM" approved="GER" date="2025-11-29" qualificationtime="00:00:33.46" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paula" lastname="Mußlick" birthdate="2006-01-01" gender="F" nation="GER" license="352742" athleteid="38201">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.27" eventid="1123" heatid="40054" lane="7">
                  <MEETINFO name="BaHaMa Cup" city="Langen" course="LCM" approved="GER" date="2025-03-22" qualificationtime="00:00:30.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.18" eventid="1207" heatid="40172" lane="8">
                  <MEETINFO name="Kreismeisterschaft Offenbach/Einlagungswettkampf" city="Heusenstamm" course="SCM" approved="GER" date="2025-11-29" qualificationtime="00:00:37.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.58" eventid="1287" heatid="40326" lane="4">
                  <MEETINFO name="BaHaMa Cup" city="Langen" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:00:31.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.58" eventid="1327" heatid="40387" lane="6">
                  <MEETINFO name="Kreismeisterschaft Offenbach/Einlagungswettkampf" city="Heusenstamm" course="SCM" approved="GER" date="2025-11-29" qualificationtime="00:01:24.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Zoé" lastname="Lempochner" birthdate="2008-01-01" gender="F" nation="GER" license="428278" athleteid="38195">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.09" eventid="1123" heatid="40039" lane="2">
                  <MEETINFO name="1. inkl. Dieburger Herbstschwimmen/13. Masters-Cup" city="Dieburg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:34.32" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.94" eventid="1143" heatid="40095" lane="4">
                  <MEETINFO name="44. Drei-Länder-Pokal" city="Lampertheim" course="SCM" approved="GER" date="2025-03-09" qualificationtime="00:03:05.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.07" eventid="1207" heatid="40170" lane="7">
                  <MEETINFO name="DMS 2024 - Bezirksliga I HSV-Süd" city="Rüsselsheim" course="SCM" approved="GER" date="2025-02-15" qualificationtime="00:00:38.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.78" eventid="1327" heatid="40388" lane="3">
                  <MEETINFO name="DMS 2024 - Bezirksliga I HSV-Süd" city="Rüsselsheim" course="SCM" approved="GER" date="2025-02-15" qualificationtime="00:01:23.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.90" eventid="1367" heatid="40447" lane="3">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:40.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Stein" birthdate="2008-01-01" gender="F" nation="GER" license="375397" athleteid="38234">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.38" eventid="1123" heatid="40044" lane="2">
                  <MEETINFO name="Bezirks- und Bezirksjahrgangsmeisterschaften" city="Darmstadt" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:00:31.38" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.02" eventid="1227" heatid="40207" lane="7">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:16.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.51" eventid="1267" heatid="40276" lane="3">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:08.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.51" eventid="1367" heatid="40452" lane="6">
                  <MEETINFO name="Bezirks- und Bezirksjahrgangsmeisterschaften" city="Darmstadt" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:35.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mara" lastname="Kutzer" birthdate="2008-01-01" gender="F" nation="GER" license="394717" athleteid="38187">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.69" eventid="1123" heatid="40042" lane="4">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:31.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.00" eventid="1163" heatid="40119" lane="3" />
                <ENTRY entrytime="00:01:21.44" eventid="1227" heatid="40201" lane="5">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:21.44" />
                </ENTRY>
                <ENTRY entrytime="00:05:00.00" eventid="1247" heatid="40243" lane="7" />
                <ENTRY entrytime="00:01:08.74" eventid="1267" heatid="40276" lane="1">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:08.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.45" eventid="1287" heatid="40315" lane="5">
                  <MEETINFO name="Bezirks- und Bezirksjahrgangsmeisterschaften" city="Darmstadt" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:00:36.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.89" eventid="1367" heatid="40445" lane="7">
                  <MEETINFO name="44. Drei-Länder-Pokal" city="Lampertheim" course="SCM" approved="GER" date="2025-03-09" qualificationtime="00:00:38.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Linda" lastname="Ogriseck" birthdate="2010-01-01" gender="F" nation="GER" license="412094" athleteid="38206">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.61" eventid="1123" heatid="40057" lane="6">
                  <MEETINFO name="Hochtaunus-Cup" city="Oberursel" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:27.61" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.76" eventid="1207" heatid="40171" lane="7">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:37.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.56" eventid="1267" heatid="40284" lane="7">
                  <MEETINFO name="Kreismeisterschaft Offenbach/Einlagungswettkampf" city="Heusenstamm" course="SCM" approved="GER" date="2025-11-29" qualificationtime="00:01:02.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.74" eventid="1287" heatid="40326" lane="3">
                  <MEETINFO name="Kreismeisterschaft Offenbach/Einlagungswettkampf" city="Heusenstamm" course="SCM" approved="GER" date="2025-11-29" qualificationtime="00:00:31.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.34" eventid="1347" heatid="40413" lane="4">
                  <MEETINFO name="Bezirks- und Bezirksjahrgangsmeisterschaften" city="Darmstadt" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:31.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Melissa" lastname="Ogriseck" birthdate="2006-01-01" gender="F" nation="GER" license="363930" athleteid="38212">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.02" eventid="1123" heatid="40057" lane="1">
                  <MEETINFO name="HM und HJM Langbahn  Darmstadt" city="Darmstadt" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:00:28.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.26" eventid="1227" heatid="40209" lane="1">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:13.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.46" eventid="1267" heatid="40284" lane="3">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:02.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.39" eventid="1287" heatid="40325" lane="6">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:31.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.55" eventid="1367" heatid="40457" lane="8">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:32.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Merle Carlotta" lastname="Knapp" birthdate="2010-01-01" gender="F" nation="GER" license="419092" athleteid="38182">
              <ENTRIES>
                <ENTRY entrytime="00:02:50.00" eventid="1143" heatid="40098" lane="4">
                  <MEETINFO name="CIJ Meet" city="Luxembourg - Kirchberg" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:03:07.75" />
                </ENTRY>
                <ENTRY entrytime="00:05:00.04" eventid="1247" heatid="40243" lane="8">
                  <MEETINFO name="1. inkl. Dieburger Herbstschwimmen/13. Masters-Cup" city="Dieburg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:05:00.04" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.85" eventid="1307" heatid="40357" lane="8">
                  <MEETINFO name="28. TSG Schwimmtest" city="Darmstadt" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:44.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.35" eventid="1347" heatid="40417" lane="7">
                  <MEETINFO name="28. TSG Schwimmtest" city="Darmstadt" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:21.97" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anastasia" lastname="Plassmann" birthdate="2009-01-01" gender="F" nation="GER" license="399719" athleteid="38218">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.24" eventid="1123" heatid="40044" lane="4">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:31.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.56" eventid="1207" heatid="40167" lane="1">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:40.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.18" eventid="1267" heatid="40272" lane="4">
                  <MEETINFO name="25. Sprintwettkampf" city="Rödermark" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:10.18" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.57" eventid="1327" heatid="40387" lane="3">
                  <MEETINFO name="DMS 2024 - Bezirksliga I HSV-Süd" city="Rüsselsheim" course="SCM" approved="GER" date="2025-02-15" qualificationtime="00:01:24.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.00" eventid="1367" heatid="40449" lane="7">
                  <MEETINFO name="BaHaMa Cup" city="Langen" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:00:39.93" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.00" eventid="1183" heatid="40144" lane="5">
                  <MEETINFO name="Kreismeisterschaft Offenbach/Einlagungswettkampf" city="Heusenstamm" date="2025-11-29" qualificationtime="00:02:15.28" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="3378" nation="GER" region="12" clubid="37876" name="SSV Leutzsch">
          <ATHLETES>
            <ATHLETE firstname="Hardy" lastname="Frank" birthdate="2011-01-01" gender="M" nation="GER" license="423159" athleteid="37890">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.42" eventid="1133" heatid="40085" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:24.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.31" eventid="1197" heatid="40154" lane="1">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:02:25.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.30" eventid="1237" heatid="40230" lane="7">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:01:03.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.16" eventid="1277" heatid="40309" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:54.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.71" eventid="1317" heatid="40374" lane="7">
                  <MEETINFO name="DMS Landesliga Berlin" city="Berlin" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:02:17.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.58" eventid="1357" heatid="40435" lane="2">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:04.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.01" eventid="1397" heatid="40494" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:00.72" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Clemens" lastname="Hartung" birthdate="2008-01-01" gender="M" nation="GER" license="368832" athleteid="37898">
              <ENTRIES>
                <ENTRY entrytime="00:02:17.86" eventid="1173" heatid="40141" lane="3">
                  <MEETINFO name="DMS Landesliga Berlin" city="Berlin" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:02:12.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.27" eventid="1197" heatid="40156" lane="2">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:02:13.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.30" eventid="1237" heatid="40231" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:00.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.21" eventid="1297" heatid="40345" lane="5">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:26.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.01" eventid="1317" heatid="40374" lane="5">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:02:23.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.86" eventid="1377" heatid="40472" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:28.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.32" eventid="1397" heatid="40496" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:58.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Richard" lastname="Plewa" birthdate="2010-01-01" gender="M" nation="GER" license="433622" athleteid="37918">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.81" eventid="1133" heatid="40084" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:26.01" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.53" eventid="1197" heatid="40153" lane="1" />
                <ENTRY entrytime="00:01:13.12" eventid="1237" heatid="40227" lane="8">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:01:14.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.71" eventid="1277" heatid="40306" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:57.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.08" eventid="1297" heatid="40344" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.73" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.35" eventid="1357" heatid="40429" lane="3" />
                <ENTRY entrytime="00:01:01.57" eventid="1397" heatid="40496" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:01.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sonja" lastname="Riemer" birthdate="2013-01-01" gender="F" nation="GER" license="461030" athleteid="37933">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.71" eventid="1123" heatid="40036" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:32.35" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.56" eventid="1163" heatid="40114" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:03:07.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.54" eventid="1207" heatid="40158" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:45.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.57" eventid="1287" heatid="40315" lane="7">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:36.57" />
                </ENTRY>
                <ENTRY entrytime="00:03:04.85" eventid="1307" heatid="40350" lane="4">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:03:04.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.06" eventid="1327" heatid="40378" lane="4">
                  <MEETINFO name="Messesprintpokal des Postschwimmverein Leipzig e.V" city="Leipzig" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:01:43.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.22" eventid="1367" heatid="40442" lane="5">
                  <MEETINFO name="Plauener Herbst- Mehrkampf" city="Plauen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:39.08" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Valentin" lastname="Plewa" birthdate="2013-01-01" gender="M" nation="GER" license="441003" athleteid="37926">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.84" eventid="1133" heatid="40073" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:29.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.38" eventid="1217" heatid="40181" lane="7">
                  <MEETINFO name="Plauener Herbst- Mehrkampf" city="Plauen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:38.38" />
                </ENTRY>
                <ENTRY entrytime="00:05:30.51" eventid="1257" heatid="40249" lane="3" />
                <ENTRY entrytime="00:01:05.13" eventid="1277" heatid="40299" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:05.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.67" eventid="1317" heatid="40369" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:38.95" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.95" eventid="1357" heatid="40428" lane="7">
                  <MEETINFO name="Giraffenpokal" city="Chemnitz" course="LCM" approved="GER" date="2025-11-08" qualificationtime="00:02:28.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Matvey" lastname="Leontyev" birthdate="2011-01-01" gender="M" nation="GER" license="418812" athleteid="37910">
              <ENTRIES>
                <ENTRY entrytime="00:02:21.51" eventid="1173" heatid="40140" lane="5">
                  <MEETINFO name="DMS Landesliga Berlin" city="Berlin" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:02:14.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.14" eventid="1197" heatid="40155" lane="7">
                  <MEETINFO name="DMS Landesliga Berlin" city="Berlin" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:02:19.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.40" eventid="1237" heatid="40230" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:02.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.60" eventid="1297" heatid="40342" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:29.60" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.50" eventid="1317" heatid="40367" lane="4" />
                <ENTRY entrytime="00:00:29.67" eventid="1377" heatid="40473" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:29.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.36" eventid="1397" heatid="40493" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:01:05.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Beyer" birthdate="2009-01-01" gender="M" nation="GER" license="382888" athleteid="37881">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.66" eventid="1133" heatid="40076" lane="4">
                  <MEETINFO name="offenes Vereinsschwimmfest" city="Eisleben" course="SCM" approved="GER" date="2025-04-26" qualificationtime="00:00:27.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.80" eventid="1173" heatid="40138" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:29.54" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.00" eventid="1197" heatid="40153" lane="6">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:02:30.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.28" eventid="1237" heatid="40229" lane="1">
                  <MEETINFO name="offenes Vereinsschwimmfest" city="Eisleben" course="SCM" approved="GER" date="2025-04-26" qualificationtime="00:01:07.38" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.76" eventid="1277" heatid="40302" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:59.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.79" eventid="1297" heatid="40342" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:29.37" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.36" eventid="1357" heatid="40431" lane="5">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:02:14.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.53" eventid="1397" heatid="40492" lane="3">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:01:05.97" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilian Arthur" lastname="Beck" birthdate="2009-01-01" gender="M" nation="GER" license="415598" athleteid="37877">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.99" eventid="1133" heatid="40086" lane="1">
                  <MEETINFO name="offenes Vereinsschwimmfest" city="Eisleben" course="SCM" approved="GER" date="2025-04-26" qualificationtime="00:00:25.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.26" eventid="1153" heatid="40107" lane="5" />
                <ENTRY entrytime="00:00:34.08" eventid="1217" heatid="40186" lane="5">
                  <MEETINFO name="Herbstschwimmfest" city="Eisleben" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:34.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Yakiv" lastname="Khrushch" birthdate="2012-01-01" gender="M" nation="GER" license="429613" athleteid="37906">
              <ENTRIES>
                <ENTRY entrytime="00:03:05.29" eventid="1153" heatid="40106" lane="1">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:03:05.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.59" eventid="1217" heatid="40180" lane="4">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:38.59" />
                </ENTRY>
                <ENTRY entrytime="00:04:43.51" eventid="1257" heatid="40256" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:04:43.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Schmidt" birthdate="2002-01-01" gender="F" nation="GER" license="263362" athleteid="37941">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.21" eventid="1123" heatid="40049" lane="1">
                  <MEETINFO name="Offene Thüringer Meisterschaften" city="Erfurt" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:30.21" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.28" eventid="1143" heatid="40096" lane="4">
                  <MEETINFO name="45. Goslarer Adler Int. Masters Schwimm Gala" city="Goslar" course="SCM" approved="GER" date="2025-03-01" qualificationtime="00:02:56.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.82" eventid="1207" heatid="40169" lane="7">
                  <MEETINFO name="Offene Thüringer Meisterschaften" city="Erfurt" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:38.82" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3351" nation="GER" region="12" clubid="38782" name="Post SV Leipzig e.V.">
          <ATHLETES>
            <ATHLETE firstname="Sanamea" lastname="Glatzel" birthdate="2008-01-01" gender="F" nation="GER" license="367036" athleteid="38783">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.88" eventid="1123" heatid="40055" lane="7">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:00:28.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.06" eventid="1143" heatid="40098" lane="6">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:02:54.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.03" eventid="1207" heatid="40173" lane="3">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:00:34.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.18" eventid="1287" heatid="40329" lane="1">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:29.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.27" eventid="1327" heatid="40390" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:01:17.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.57" eventid="1367" heatid="40456" lane="4">
                  <MEETINFO name="44.Wettbewerb um die Mehrkampfpokale" city="Leipzig" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:33.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4949" nation="GER" region="07" clubid="35811" name="SG Wetterau">
          <ATHLETES>
            <ATHLETE firstname="Lukas" lastname="Margraf" birthdate="2012-01-01" gender="M" nation="GER" license="453756" athleteid="35818">
              <ENTRIES>
                <ENTRY entrytime="00:09:33.01" eventid="1093" heatid="40018" lane="1">
                  <MEETINFO name="Hochtaunus-Cup" city="Oberursel" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:09:33.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.35" eventid="1133" heatid="40078" lane="2">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:28.35" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.36" eventid="1173" heatid="40137" lane="2">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:02:39.66" />
                </ENTRY>
                <ENTRY entrytime="00:04:39.86" eventid="1257" heatid="40258" lane="8">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:04:39.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.07" eventid="1277" heatid="40302" lane="8">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:03.07" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.99" eventid="1357" heatid="40433" lane="4">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:02:13.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Victoria Louise" lastname="Humann" birthdate="2015-01-01" gender="F" nation="GER" license="467709" athleteid="35812">
              <ENTRIES>
                <ENTRY entrytime="00:03:14.27" eventid="1143" heatid="40093" lane="4">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:03:14.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.41" eventid="1207" heatid="40159" lane="8">
                  <MEETINFO name="HM und HJM Langbahn  Darmstadt" city="Darmstadt" course="LCM" approved="GER" date="2025-06-20" qualificationtime="00:00:45.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.58" eventid="1287" heatid="40313" lane="1">
                  <MEETINFO name="Bezirksmeisterschaft - HSV Bezirk Mitte" city="Offenbach" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:00:39.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.04" eventid="1327" heatid="40381" lane="2">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:34.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.55" eventid="1387" heatid="40477" lane="7">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:30.55" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Justus Florian" lastname="Rose" birthdate="2007-01-01" gender="M" nation="GER" license="387915" athleteid="35825">
              <ENTRIES>
                <ENTRY entrytime="00:02:35.91" eventid="1153" heatid="40110" lane="3">
                  <MEETINFO name="37. Herbstpokal der SG Frankfurt" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:02:35.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.59" eventid="1217" heatid="40188" lane="4">
                  <MEETINFO name="Internationales Frühjahrsmeeting SG Wetterau" city="Bad Nauheim" course="LCM" approved="GER" date="2025-05-01" qualificationtime="00:00:31.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.17" eventid="1277" heatid="40308" lane="3">
                  <MEETINFO name="Hochtaunus-Cup" city="Oberursel" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:58.17" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.99" eventid="1337" heatid="40402" lane="2">
                  <MEETINFO name="HM und HJM Langbahn  Darmstadt" city="Darmstadt" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:10.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Salome" lastname="Schultheis" birthdate="2008-01-01" gender="F" nation="GER" license="379210" athleteid="35830">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.38" eventid="1123" heatid="40049" lane="8">
                  <MEETINFO name="BaHaMa Cup" city="Langen" course="LCM" approved="GER" date="2025-03-22" qualificationtime="00:00:30.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.28" eventid="1207" heatid="40168" lane="7">
                  <MEETINFO name="Hochtaunus-Cup" city="Oberursel" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:39.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.78" eventid="1287" heatid="40326" lane="2">
                  <MEETINFO name="Bezirksmeisterschaft - HSV Bezirk Mitte" city="Offenbach" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:00:31.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.91" eventid="1387" heatid="40483" lane="8">
                  <MEETINFO name="HM und HJM Langbahn  Darmstadt" city="Darmstadt" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:13.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Trautmann" birthdate="2009-01-01" gender="F" nation="GER" license="443502" athleteid="35835">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.55" eventid="1123" heatid="40048" lane="7">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:30.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.51" eventid="1163" heatid="40121" lane="1">
                  <MEETINFO name="37. Herbstpokal der SG Frankfurt" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:02:47.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.24" eventid="1227" heatid="40206" lane="8">
                  <MEETINFO name="Hochtaunus-Cup" city="Oberursel" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:17.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.93" eventid="1267" heatid="40273" lane="6">
                  <MEETINFO name="BaHaMa Cup" city="Langen" course="LCM" approved="GER" date="2025-03-22" qualificationtime="00:01:09.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.37" eventid="1367" heatid="40454" lane="4">
                  <MEETINFO name="HM und HJM Kurzbahn  Fulda" city="Fulda" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:34.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Ramona" gender="M" lastname="Kerkhoff" />
            <COACH firstname="Stefan" gender="M" lastname="Kaul" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="00000" nation="AUT" clubid="38141" name="Tiroler Wassersportverein">
          <ATHLETES>
            <ATHLETE firstname="Rosa" lastname="Maier-Dejaco" birthdate="2011-01-01" gender="F" nation="AUT" license="0" athleteid="38151">
              <ENTRIES>
                <ENTRY entrytime="00:03:13.50" eventid="1143" heatid="40094" lane="8" />
                <ENTRY entrytime="00:00:39.98" eventid="1207" heatid="40166" lane="5" />
                <ENTRY entrytime="00:01:25.48" eventid="1227" heatid="40197" lane="7" />
                <ENTRY entrytime="00:01:14.38" eventid="1267" heatid="40267" lane="3" />
                <ENTRY entrytime="00:01:30.06" eventid="1327" heatid="40383" lane="6" />
                <ENTRY entrytime="00:00:41.73" eventid="1367" heatid="40441" lane="3" />
                <ENTRY entrytime="00:01:24.73" eventid="1387" heatid="40478" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Kim" lastname="Koller" birthdate="2010-01-01" gender="F" nation="AUT" license="0" athleteid="38159">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.84" eventid="1123" heatid="40047" lane="8" />
                <ENTRY entrytime="00:02:49.23" eventid="1163" heatid="40120" lane="2" />
                <ENTRY entrytime="00:01:18.20" eventid="1227" heatid="40205" lane="1" />
                <ENTRY entrytime="00:01:11.12" eventid="1267" heatid="40271" lane="3" />
                <ENTRY entrytime="00:00:33.93" eventid="1287" heatid="40321" lane="7" />
                <ENTRY entrytime="00:00:36.43" eventid="1367" heatid="40450" lane="6" />
                <ENTRY entrytime="00:01:17.85" eventid="1387" heatid="40480" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Blaukovitsch" birthdate="2010-01-01" gender="F" nation="AUT" license="0" athleteid="38167">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.12" eventid="1123" heatid="40035" lane="7" />
                <ENTRY entrytime="00:00:41.76" eventid="1207" heatid="40163" lane="4" />
                <ENTRY entrytime="00:01:13.38" eventid="1267" heatid="40268" lane="5" />
                <ENTRY entrytime="00:01:35.96" eventid="1327" heatid="40380" lane="3" />
                <ENTRY entrytime="00:02:46.41" eventid="1347" heatid="40407" lane="4" />
                <ENTRY entrytime="00:00:42.87" eventid="1367" heatid="40440" lane="5" />
                <ENTRY entrytime="00:00:41.52" eventid="1287" heatid="40312" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Eichholzer" birthdate="2007-01-01" gender="F" nation="AUT" license="0" athleteid="38142">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.27" eventid="1123" heatid="40054" lane="1" />
                <ENTRY entrytime="00:03:05.67" eventid="1143" heatid="40096" lane="1" />
                <ENTRY entrytime="00:00:40.00" eventid="1207" heatid="40166" lane="3" />
                <ENTRY entrytime="00:01:19.32" eventid="1227" heatid="40204" lane="2" />
                <ENTRY entrytime="00:01:06.05" eventid="1267" heatid="40279" lane="3" />
                <ENTRY entrytime="00:00:31.32" eventid="1287" heatid="40327" lane="6" />
                <ENTRY entrytime="00:02:26.59" eventid="1347" heatid="40416" lane="1" />
                <ENTRY entrytime="00:01:18.86" eventid="1387" heatid="40480" lane="8" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1183" heatid="40143" lane="2" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="3580" nation="GER" region="13" clubid="38544" name="SC Magdeburg">
          <ATHLETES>
            <ATHLETE firstname="Maximilian" lastname="Kraus" birthdate="2014-01-01" gender="M" nation="GER" license="443519" athleteid="38570">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.07" eventid="1133" heatid="40070" lane="4">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:31.07" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.43" eventid="1173" heatid="40135" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:45.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.46" eventid="1237" heatid="40224" lane="8">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:01:17.46" />
                </ENTRY>
                <ENTRY entrytime="00:05:06.03" eventid="1257" heatid="40253" lane="4">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:05:04.21" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.81" eventid="1277" heatid="40297" lane="5">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:01:07.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.94" eventid="1297" heatid="40335" lane="4">
                  <MEETINFO name="Kids-Cup Teil 1 des LSVSA der Leistungsstützpunkte" city="Bitterfeld-Wolfen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:34.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Laia" lastname="Gutiérrez Müller" birthdate="2012-01-01" gender="F" nation="GER" license="476631" athleteid="38560">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.90" eventid="1287" status="WDR">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:30.90" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.55" eventid="1327" status="WDR">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:21.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.00" eventid="1347" status="WDR">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:20.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.33" eventid="1367" status="WDR">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:33.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lotta" lastname="Adam" birthdate="2010-01-01" gender="F" nation="GER" license="414440" athleteid="38545">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.30" eventid="1267" heatid="40284" lane="5">
                  <MEETINFO name="DMSJ" city="Burg" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:00.14" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.45" eventid="1327" heatid="40386" lane="5">
                  <MEETINFO name="DMSJ" city="Burg" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:19.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.01" eventid="1367" heatid="40459" lane="6">
                  <MEETINFO name="Lagen - Wettkampf" city="Magdeburg" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:00:32.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.54" eventid="1387" heatid="40484" lane="5">
                  <MEETINFO name="DMSJ" city="Burg" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:07.82" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marlene" lastname="Himmel" birthdate="2011-01-01" gender="F" nation="GER" license="442520" athleteid="38565">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.55" eventid="1287" heatid="40317" lane="7">
                  <MEETINFO name="34. Gothaer &amp; Friends mit Kids Pokal" city="Magdeburg" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:00:35.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.28" eventid="1327" heatid="40385" lane="5">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:01:31.99" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.48" eventid="1347" heatid="40416" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:24.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.82" eventid="1367" heatid="40456" lane="7">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:32.87" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Constantin" lastname="Fabian" birthdate="2011-01-01" gender="M" nation="GER" license="430675" athleteid="38555">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.30" eventid="1277" heatid="40305" lane="3">
                  <MEETINFO name="DMSJ" city="Burg" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:57.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.90" eventid="1337" heatid="40400" lane="4">
                  <MEETINFO name="DMSJ" city="Burg" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:10.35" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.62" eventid="1357" heatid="40433" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:14.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.33" eventid="1377" heatid="40471" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Eva" lastname="Woitag" birthdate="2011-01-01" gender="F" nation="GER" license="387151" athleteid="38607">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.50" eventid="1287" heatid="40329" lane="3">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:00:27.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.40" eventid="1327" heatid="40388" lane="4">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:23.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.72" eventid="1347" heatid="40420" lane="2">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:02:04.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.21" eventid="1367" heatid="40459" lane="4">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:30.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maximilian" lastname="Wiemer" birthdate="2010-01-01" gender="M" nation="GER" license="409856" athleteid="38602">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.58" eventid="1277" heatid="40310" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:56.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.55" eventid="1337" heatid="40401" lane="1">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:16.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.89" eventid="1357" heatid="40437" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:05.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.12" eventid="1377" heatid="40472" lane="1">
                  <MEETINFO name="Lagen - Wettkampf" city="Magdeburg" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:00:31.12" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Katharina" lastname="Slach" birthdate="2012-01-01" gender="F" nation="GER" license="436752" athleteid="38592">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.15" eventid="1267" heatid="40279" lane="8">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:01:07.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.62" eventid="1287" heatid="40321" lane="5">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:33.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.21" eventid="1347" heatid="40417" lane="1">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:24.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.33" eventid="1367" heatid="40450" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lisa" lastname="Barth" birthdate="2010-01-01" gender="F" nation="GER" license="377094" athleteid="38550">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.04" eventid="1267" heatid="40286" lane="7">
                  <MEETINFO name="34. Gothaer &amp; Friends mit Kids Pokal" city="Magdeburg" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:01:00.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.77" eventid="1327" heatid="40389" lane="3" />
                <ENTRY entrytime="00:02:11.03" eventid="1347" heatid="40420" lane="8">
                  <MEETINFO name="Überprüfungswettkampf" city="Halle (Saale)" course="LCM" approved="GER" date="2025-02-08" qualificationtime="00:02:11.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.79" eventid="1367" heatid="40457" lane="5">
                  <MEETINFO name="Lagen - Wettkampf" city="Magdeburg" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:00:32.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Schmidt" birthdate="2010-01-01" gender="M" nation="GER" license="409854" athleteid="38587">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.20" eventid="1277" heatid="40307" lane="2">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:01:02.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.07" eventid="1297" heatid="40343" lane="7">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:00:29.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.95" eventid="1337" heatid="40401" lane="3">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:12.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.10" eventid="1357" heatid="40433" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:14.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Laura Eszter" lastname="Toth" birthdate="2012-01-01" gender="F" nation="GER" license="436388" athleteid="38597">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.03" eventid="1267" heatid="40282" lane="6">
                  <MEETINFO name="34. Gothaer &amp; Friends mit Kids Pokal" city="Magdeburg" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:01:04.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.33" eventid="1327" heatid="40386" lane="6" />
                <ENTRY entrytime="00:02:19.09" eventid="1347" heatid="40418" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:19.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.75" eventid="1367" heatid="40454" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mattis" lastname="Nebelung" birthdate="2009-01-01" gender="M" nation="GER" license="369734" athleteid="38582">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.16" eventid="1277" heatid="40308" lane="5">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:56.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.65" eventid="1297" heatid="40343" lane="4">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:27.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.41" eventid="1357" heatid="40436" lane="7">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:02:03.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.18" eventid="1377" heatid="40473" lane="2">
                  <MEETINFO name="35. Dompfaff-Pokal Fulda" city="Fulda" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:28.97" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Artemiy" lastname="Kuzmin" birthdate="2011-01-01" gender="M" nation="GER" license="426385" athleteid="38577">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.05" eventid="1297" heatid="40339" lane="1">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:32.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.08" eventid="1337" heatid="40399" lane="3">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:01:19.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.66" eventid="1357" heatid="40430" lane="4">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:20.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.49" eventid="1377" heatid="40466" lane="8" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4738" nation="GER" region="04" clubid="35903" name="SSV PCK 90 Schwedt">
          <ATHLETES>
            <ATHLETE firstname="Marie" lastname="Lienert" birthdate="2011-01-01" gender="F" nation="GER" license="423581" athleteid="35926">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.68" eventid="1123" heatid="40033" lane="2">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:33.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.04" eventid="1207" heatid="40162" lane="4">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:42.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.36" eventid="1267" heatid="40266" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:15.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.56" eventid="1287" heatid="40315" lane="2">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:00:36.56" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Cedric" lastname="Sasse" birthdate="2008-01-01" gender="M" nation="GER" license="379485" athleteid="35949">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.62" eventid="1133" heatid="40084" lane="6">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:26.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.35" eventid="1217" heatid="40188" lane="2">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:31.50" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.08" eventid="1317" heatid="40374" lane="3" />
                <ENTRY entrytime="00:01:12.16" eventid="1337" heatid="40402" lane="1">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:09.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nela" lastname="Willim" birthdate="2013-01-01" gender="F" nation="GER" license="446938" athleteid="35971">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.55" eventid="1123" heatid="40031" lane="2">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:32.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.46" eventid="1227" heatid="40195" lane="8">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:22.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.31" eventid="1267" heatid="40264" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:13.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.79" eventid="1287" heatid="40314" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:36.79" />
                </ENTRY>
                <ENTRY entrytime="00:03:11.68" eventid="1307" heatid="40349" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:03:04.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.25" eventid="1367" heatid="40444" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:39.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sarah-Sophie" lastname="Matern" birthdate="2008-01-01" gender="F" nation="GER" license="379495" athleteid="35938">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.39" eventid="1123" heatid="40037" lane="6">
                  <MEETINFO name="26. Int. Berolina Cup" city="Berlin" course="LCM" approved="GER" date="2025-02-22" qualificationtime="00:00:32.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.79" eventid="1267" heatid="40270" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:11.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.41" eventid="1287" heatid="40315" lane="4">
                  <MEETINFO name="26. Int. Berolina Cup" city="Berlin" course="LCM" approved="GER" date="2025-02-23" qualificationtime="00:00:36.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Tabea" lastname="Sasse" birthdate="2004-01-01" gender="F" nation="GER" license="315166" athleteid="35954">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.75" eventid="1123" heatid="40047" lane="1">
                  <MEETINFO name="Offene Berliner Kurzbahnmeisterschaften Masters" city="Berlin" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:00:30.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.77" eventid="1207" heatid="40172" lane="2">
                  <MEETINFO name="Offene Berliner Kurzbahnmeisterschaften Masters" city="Berlin" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:00:36.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.15" eventid="1287" heatid="40327" lane="3">
                  <MEETINFO name="Offene Berliner Kurzbahnmeisterschaften Masters" city="Berlin" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:00:31.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.36" eventid="1327" heatid="40388" lane="8">
                  <MEETINFO name="XIX. Rostock Masters Sprint Cup" city="Rostock" course="SCM" approved="GER" date="2025-06-21" qualificationtime="00:01:21.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Tinginies" birthdate="2013-01-01" gender="F" nation="GER" license="447021" athleteid="35959">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.84" eventid="1123" heatid="40036" lane="7">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:32.03" />
                </ENTRY>
                <ENTRY entrytime="00:03:35.64" eventid="1143" heatid="40090" lane="5">
                  <MEETINFO name="16. Internationales Nachwuchsschwimmfest" city="Cottbus" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:03:35.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.83" eventid="1207" heatid="40159" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:42.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.44" eventid="1227" heatid="40196" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:24.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.05" eventid="1267" heatid="40270" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:12.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.63" eventid="1327" heatid="40380" lane="2">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:34.47" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.77" eventid="1347" heatid="40407" lane="3">
                  <MEETINFO name="Barnim-Uckermark Cup" city="Eberswalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:48.77" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="John" lastname="Lienert" birthdate="2008-01-01" gender="M" nation="GER" license="379486" athleteid="35921">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.80" eventid="1133" heatid="40074" lane="1">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:00:29.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.63" eventid="1277" heatid="40298" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:06.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.11" eventid="1297" heatid="40340" lane="8">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:00:31.11" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.94" eventid="1397" heatid="40491" lane="6">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:10.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Otto" birthdate="2002-01-01" gender="F" nation="GER" license="300972" athleteid="35942">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.83" eventid="1123" heatid="40041" lane="3">
                  <MEETINFO name="Offene Berliner Kurzbahnmeisterschaften Masters" city="Berlin" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:00:32.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Victoria" lastname="Putzke" birthdate="2010-01-01" gender="F" nation="GER" license="414209" athleteid="35944">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.13" eventid="1123" heatid="40050" lane="8">
                  <MEETINFO name="Barnim-Uckermark Cup" city="Eberswalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:00:29.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.87" eventid="1207" heatid="40169" lane="1">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:38.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.57" eventid="1287" heatid="40324" lane="5">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:00:32.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.14" eventid="1327" heatid="40389" lane="8">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:23.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Malea" lastname="Willim" birthdate="2008-01-01" gender="F" nation="GER" license="379488" athleteid="35967">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.99" eventid="1123" heatid="40032" lane="6">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:33.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.89" eventid="1207" heatid="40165" lane="7">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:40.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.96" eventid="1327" heatid="40383" lane="3">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:29.96" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Stella-Lotte" lastname="Krauße" birthdate="2011-01-01" gender="F" nation="GER" license="436568" athleteid="35916">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.72" eventid="1123" heatid="40033" lane="7">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:33.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.70" eventid="1207" heatid="40160" lane="8">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:44.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.35" eventid="1267" heatid="40267" lane="5">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:14.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.90" eventid="1327" heatid="40382" lane="1">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:31.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Luna Victoria" lastname="Fatke" birthdate="2013-01-01" gender="F" nation="GER" license="446917" athleteid="35904">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.49" eventid="1123" heatid="40034" lane="1">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:32.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.11" eventid="1227" heatid="40198" lane="5">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:21.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.00" eventid="1267" heatid="40269" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:11.52" />
                </ENTRY>
                <ENTRY entrytime="00:03:08.70" eventid="1307" heatid="40349" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:03:05.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.63" eventid="1367" heatid="40445" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:37.82" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Janis" lastname="Lück" birthdate="2013-01-01" gender="M" nation="GER" license="446940" athleteid="35931">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.25" eventid="1133" heatid="40066" lane="7">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:31.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.13" eventid="1237" heatid="40220" lane="3" />
                <ENTRY entrytime="00:01:11.32" eventid="1277" heatid="40295" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:09.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.37" eventid="1297" heatid="40337" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:33.37" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.63" eventid="1317" heatid="40369" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:45.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.59" eventid="1377" heatid="40467" lane="1">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:35.46" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jonas" lastname="Kleinke" birthdate="2008-01-01" gender="M" nation="GER" license="386677" athleteid="35910">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.82" eventid="1133" heatid="40080" lane="1">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:27.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.19" eventid="1173" heatid="40138" lane="7" />
                <ENTRY entrytime="00:01:09.16" eventid="1237" heatid="40229" lane="5">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:06.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.00" eventid="1277" heatid="40302" lane="6">
                  <MEETINFO name="Forstpokal" city="Eberswalde" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:59.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.24" eventid="1377" heatid="40471" lane="5">
                  <MEETINFO name="MV-Cup Vorkampf in Neubrandenburg" city="Neubrandenburg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:30.80" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Lea" gender="M" lastname="Otto" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="5129" nation="GER" region="14" clubid="34932" name="SV Neptun Kiel">
          <ATHLETES>
            <ATHLETE firstname="Finn-Luca" lastname="Malcherek" birthdate="2013-01-01" gender="M" nation="GER" license="446591" athleteid="34984">
              <ENTRIES>
                <ENTRY entrytime="00:10:40.00" eventid="1093" heatid="40014" lane="4" />
                <ENTRY entrytime="00:00:34.46" eventid="1133" heatid="40064" lane="1">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:34.34" />
                </ENTRY>
                <ENTRY entrytime="00:03:29.10" eventid="1153" heatid="40103" lane="8">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:03:25.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.53" eventid="1217" heatid="40178" lane="6">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:42.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.50" eventid="1277" heatid="40290" lane="1">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:01:16.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.13" eventid="1337" heatid="40393" lane="2">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:01:37.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.67" eventid="1357" heatid="40422" lane="7">
                  <MEETINFO name="1. Swim-Cup powered by Stadtwerke Solingen" city="Solingen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:58.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.59" eventid="1377" heatid="40461" lane="7">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:42.12" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Swana" lastname="Stawczynski" birthdate="2015-01-01" gender="F" nation="GER" license="455881" athleteid="35035">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.63" eventid="1123" heatid="40026" lane="3">
                  <MEETINFO name="SHSV-Sprintmehrkampf &amp; Staffel-MS" city="Lübeck" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:38.23" />
                </ENTRY>
                <ENTRY entrytime="00:03:44.00" eventid="1163" heatid="40112" lane="7">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:03:44.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.98" eventid="1207" heatid="40157" lane="6">
                  <MEETINFO name="SHSV-Sprintmehrkampf &amp; Staffel-MS" city="Lübeck" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:54.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.26" eventid="1227" heatid="40191" lane="5">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:42.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.55" eventid="1267" heatid="40262" lane="7">
                  <MEETINFO name="SHSV-MS, JG-MS und SMK" city="Kiel" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:01:23.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.14" eventid="1327" heatid="40377" lane="3">
                  <MEETINFO name="DMS-J Landesentscheid" city="Niebüll" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:01.72" />
                </ENTRY>
                <ENTRY entrytime="00:03:04.74" eventid="1347" heatid="40405" lane="1">
                  <MEETINFO name="SHSV-MS, JG-MS und SMK" city="Kiel" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:03:04.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.20" eventid="1367" heatid="40439" lane="3">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:00:47.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lotta" lastname="Göttsche" birthdate="2002-01-01" gender="F" nation="GER" license="302745" athleteid="34951">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.29" eventid="1123" heatid="40056" lane="2">
                  <MEETINFO name="32. Sommerwettkämpfe mit dem 1. Kieler-Woche-Pokal" city="Kiel" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:27.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.96" eventid="1163" heatid="40124" lane="4">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:30.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.25" eventid="1227" heatid="40211" lane="1">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:07.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.17" eventid="1267" heatid="40282" lane="1">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:01.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.95" eventid="1367" heatid="40459" lane="8">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:31.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hanne" lastname="Wigger" birthdate="2009-01-01" gender="F" nation="GER" license="436425" athleteid="35075">
              <ENTRIES>
                <ENTRY entrytime="00:10:00.50" eventid="1083" heatid="40011" lane="8" />
                <ENTRY entrytime="00:00:29.28" eventid="1123" heatid="40054" lane="8">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:29.28" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.18" eventid="1163" heatid="40122" lane="3">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:43.18" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.82" eventid="1227" heatid="40207" lane="6">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:15.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.17" eventid="1267" heatid="40282" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:04.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.50" eventid="1287" heatid="40324" lane="4">
                  <MEETINFO name="Bille Cup" city="Lübeck" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:33.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.40" eventid="1367" heatid="40450" lane="3">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:35.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emma Sophie" lastname="Domm" birthdate="2014-01-01" gender="F" nation="GER" license="455486" athleteid="34933">
              <ENTRIES>
                <ENTRY entrytime="00:11:45.99" eventid="1083" heatid="40004" lane="7">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:11:21.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.72" eventid="1123" heatid="40029" lane="8">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:32.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.38" eventid="1163" heatid="40118" lane="6">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:02:53.38" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.81" eventid="1227" heatid="40193" lane="3">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:01:20.70" />
                </ENTRY>
                <ENTRY entrytime="00:05:36.86" eventid="1247" heatid="40237" lane="1">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:05:26.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.75" eventid="1267" heatid="40266" lane="3">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:11.76" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.35" eventid="1307" heatid="40350" lane="1">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:03:03.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.81" eventid="1347" heatid="40408" lane="3">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:02:33.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.15" eventid="1367" heatid="40441" lane="4">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:38.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ella" lastname="Weber" birthdate="2013-01-01" gender="F" nation="GER" license="473789" athleteid="35057">
              <ENTRIES>
                <ENTRY entrytime="00:21:30.00" eventid="1103" heatid="40021" lane="1" />
                <ENTRY entrytime="00:00:33.45" eventid="1123" heatid="40034" lane="2">
                  <MEETINFO name="SHSV-Sprintmehrkampf &amp; Staffel-MS" city="Lübeck" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:33.38" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.85" eventid="1163" heatid="40117" lane="2">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:47.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.62" eventid="1227" heatid="40198" lane="7">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:19.17" />
                </ENTRY>
                <ENTRY entrytime="00:05:22.37" eventid="1247" heatid="40238" lane="5">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:05:12.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.09" eventid="1267" heatid="40268" lane="4">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:09.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.46" eventid="1307" heatid="40354" lane="1">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:49.75" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.02" eventid="1347" heatid="40411" lane="3">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:30.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.37" eventid="1367" heatid="40444" lane="7">
                  <MEETINFO name="SHSV-Sprintmehrkampf &amp; Staffel-MS" city="Lübeck" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:38.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Silas" lastname="Quickert" birthdate="2014-01-01" gender="M" nation="GER" license="455489" athleteid="34993">
              <ENTRIES>
                <ENTRY entrytime="00:11:10.00" eventid="1093" heatid="40013" lane="4" />
                <ENTRY entrytime="00:00:33.42" eventid="1133" heatid="40065" lane="5">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:30.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.88" eventid="1173" heatid="40133" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:54.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.40" eventid="1217" heatid="40175" lane="5">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:41.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.17" eventid="1237" heatid="40216" lane="3">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:19.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.09" eventid="1277" heatid="40292" lane="8">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:10.71" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.73" eventid="1337" heatid="40391" lane="3">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:32.77" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.53" eventid="1357" heatid="40423" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:32.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.80" eventid="1377" heatid="40463" lane="3">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:37.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Bo Bent Arvid" lastname="Hecker" birthdate="2007-01-01" gender="M" nation="GER" license="389660" athleteid="34957">
              <ENTRIES>
                <ENTRY entrytime="00:10:51.12" eventid="1093" heatid="40014" lane="7">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:09:55.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.23" eventid="1133" heatid="40075" lane="3">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:27.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.82" eventid="1217" heatid="40180" lane="3" />
                <ENTRY entrytime="00:01:20.05" eventid="1237" heatid="40222" lane="7" />
                <ENTRY entrytime="00:06:28.68" eventid="1257" heatid="40246" lane="6" />
                <ENTRY entrytime="00:01:04.96" eventid="1277" heatid="40299" lane="4" />
                <ENTRY entrytime="00:02:24.46" eventid="1357" heatid="40429" lane="6">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:14.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.32" eventid="1377" heatid="40466" lane="1">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:33.68" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Frieda" lastname="Voss" birthdate="2011-01-01" gender="F" nation="GER" license="433402" athleteid="35050">
              <ENTRIES>
                <ENTRY entrytime="00:11:38.22" eventid="1083" heatid="40004" lane="3" />
                <ENTRY entrytime="00:00:29.26" eventid="1123" heatid="40054" lane="2">
                  <MEETINFO name="32. Sommerwettkämpfe mit dem 1. Kieler-Woche-Pokal" city="Kiel" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:28.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.72" eventid="1227" heatid="40200" lane="2">
                  <MEETINFO name="32. Winterwettkämpfe" city="Kiel" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:01:22.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.81" eventid="1267" heatid="40280" lane="8">
                  <MEETINFO name="32. Sommerwettkämpfe mit dem 1. Kieler-Woche-Pokal" city="Kiel" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:05.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.70" eventid="1287" heatid="40328" lane="4">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:29.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.32" eventid="1387" heatid="40482" lane="1">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:09.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karolin" lastname="Schlotfeldt" birthdate="2012-01-01" gender="F" nation="GER" license="474837" athleteid="35021">
              <ENTRIES>
                <ENTRY entrytime="00:11:27.50" eventid="1083" heatid="40005" lane="3" />
                <ENTRY entrytime="00:00:30.65" eventid="1123" heatid="40047" lane="5">
                  <MEETINFO name="SHSV-Sprintmehrkampf &amp; Staffel-MS" city="Lübeck" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:30.65" />
                </ENTRY>
                <ENTRY entrytime="00:03:15.34" eventid="1143" heatid="40093" lane="5">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:03:05.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.57" eventid="1207" heatid="40166" lane="8">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:40.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.75" eventid="1267" heatid="40277" lane="5">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:07.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.85" eventid="1287" heatid="40318" lane="3">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:33.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.00" eventid="1327" heatid="40384" lane="2">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:28.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.52" eventid="1387" heatid="40482" lane="8">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:13.98" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Tino" lastname="Riecken" birthdate="2012-01-01" gender="M" nation="GER" license="442207" athleteid="35003">
              <ENTRIES>
                <ENTRY entrytime="00:10:30.00" eventid="1093" heatid="40015" lane="6" />
                <ENTRY entrytime="00:00:30.77" eventid="1133" heatid="40071" lane="6">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:28.86" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.45" eventid="1153" heatid="40105" lane="6">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:55.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.18" eventid="1217" heatid="40182" lane="5">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:00:35.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.29" eventid="1317" heatid="40367" lane="3">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:39.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.59" eventid="1337" heatid="40397" lane="8">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:17.72" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.82" eventid="1357" heatid="40426" lane="1">
                  <MEETINFO name="Neptun Schwimmfest" city="Kiel" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:02:35.82" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lotta Marie" lastname="Stratmann" birthdate="2009-01-01" gender="F" nation="GER" license="398686" athleteid="35044">
              <ENTRIES>
                <ENTRY entrytime="00:10:15.30" eventid="1083" heatid="40010" lane="8" />
                <ENTRY entrytime="00:00:30.15" eventid="1123" heatid="40049" lane="5">
                  <MEETINFO name="SHSV-MS, JG-MS und SMK" city="Kiel" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:00:30.48" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.84" eventid="1187" heatid="40150" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:43.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.89" eventid="1287" heatid="40328" lane="6">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:30.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.71" eventid="1387" heatid="40484" lane="3">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:08.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emma Sophie" lastname="Wright" birthdate="2009-01-01" gender="F" nation="GER" license="442601" athleteid="35083">
              <ENTRIES>
                <ENTRY entrytime="00:10:10.00" eventid="1083" heatid="40010" lane="2" />
                <ENTRY entrytime="00:00:34.14" eventid="1123" heatid="40032" lane="7">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:31.99" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.98" eventid="1163" heatid="40121" lane="6">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:45.98" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.89" eventid="1227" heatid="40206" lane="2">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:16.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.37" eventid="1267" heatid="40274" lane="2">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:01:09.37" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.46" eventid="1287" heatid="40319" lane="6">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:00:34.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.57" eventid="1367" heatid="40450" lane="8">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:00:36.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.88" eventid="1387" heatid="40479" lane="4">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:18.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Amelie" lastname="Rother" birthdate="2014-01-01" gender="F" nation="GER" license="473316" athleteid="35011">
              <ENTRIES>
                <ENTRY entrytime="00:11:35.00" eventid="1083" heatid="40004" lane="4">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:12:44.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.42" eventid="1123" heatid="40029" lane="6">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:32.99" />
                </ENTRY>
                <ENTRY entrytime="00:03:09.31" eventid="1143" heatid="40094" lane="4">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:03:09.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.91" eventid="1207" heatid="40167" lane="8">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:38.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.76" eventid="1227" heatid="40200" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:22.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.38" eventid="1267" heatid="40265" lane="1">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:16.71" />
                </ENTRY>
                <ENTRY entrytime="00:03:18.08" eventid="1307" heatid="40349" lane="1">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:03:02.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.14" eventid="1327" heatid="40385" lane="8">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:26.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.50" eventid="1347" heatid="40407" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Holly Marie" lastname="Weinke" birthdate="2007-01-01" gender="F" nation="GER" license="358378" athleteid="35067">
              <ENTRIES>
                <ENTRY entrytime="00:09:50.00" eventid="1083" heatid="40011" lane="7" />
                <ENTRY entrytime="00:02:59.41" eventid="1163" heatid="40116" lane="2">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:02:59.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.86" eventid="1207" heatid="40161" lane="5">
                  <MEETINFO name="32. Wiking-Pokal" city="Kiel" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:47.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.64" eventid="1227" heatid="40198" lane="1">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:24.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.50" eventid="1287" heatid="40319" lane="1">
                  <MEETINFO name="32. Wiking-Pokal" city="Kiel" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:40.38" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.34" eventid="1307" heatid="40350" lane="7" />
                <ENTRY entrytime="00:00:38.15" eventid="1367" heatid="40446" lane="4">
                  <MEETINFO name="32. Wiking-Pokal" city="Kiel" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:39.12" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hans Mathis" lastname="Sommer" birthdate="2004-01-01" gender="M" nation="GER" license="324659" athleteid="35030">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.91" eventid="1133" heatid="40086" lane="6">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:26.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.94" eventid="1217" heatid="40188" lane="6">
                  <MEETINFO name="SHSV-MS, JG-MS und SMK" city="Kiel" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:00:32.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.76" eventid="1297" heatid="40346" lane="5">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:26.37" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.40" eventid="1397" heatid="40496" lane="1">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:00.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Phibie-Frederike" lastname="Dücker" birthdate="2008-01-01" gender="F" nation="GER" license="386729" athleteid="34943">
              <ENTRIES>
                <ENTRY entrytime="00:05:31.41" eventid="1063" heatid="39996" lane="4">
                  <MEETINFO name="Norddeutsche Meisterschaften Lange Strecken" city="Braunschweig" course="LCM" approved="GER" date="2025-02-15" qualificationtime="00:05:33.82" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.38" eventid="1123" heatid="40056" lane="1">
                  <MEETINFO name="32. Sommerwettkämpfe mit dem 1. Kieler-Woche-Pokal" city="Kiel" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:28.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.79" eventid="1163" heatid="40124" lane="2">
                  <MEETINFO name="32. Winterwettkämpfe" city="Kiel" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:02:45.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.00" eventid="1207" heatid="40172" lane="3">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:35.14" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.75" eventid="1267" heatid="40284" lane="4">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:02.34" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.20" eventid="1307" heatid="40360" lane="2">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:27.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.40" eventid="1347" heatid="40419" lane="1">
                  <MEETINFO name="32. Winterwettkämpfe" city="Kiel" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:02:19.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Levke" lastname="Krüger" birthdate="2008-01-01" gender="F" nation="GER" license="397492" athleteid="34966">
              <ENTRIES>
                <ENTRY entrytime="00:19:23.21" eventid="1103" heatid="40021" lane="3">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:19:12.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.89" eventid="1123" heatid="40050" lane="4" />
                <ENTRY entrytime="00:02:32.82" eventid="1163" heatid="40126" lane="1">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:02:29.22" />
                </ENTRY>
                <ENTRY entrytime="00:04:54.25" eventid="1247" heatid="40243" lane="5">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:04:43.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.25" eventid="1267" heatid="40282" lane="8">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:03.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.84" eventid="1347" heatid="40418" lane="6">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:15.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.58" eventid="1367" heatid="40456" lane="5">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:33.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Rieke" lastname="Krüger" birthdate="2012-01-01" gender="F" nation="GER" license="408719" athleteid="34974">
              <ENTRIES>
                <ENTRY entrytime="00:11:01.76" eventid="1083" heatid="40007" lane="8">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:10:23.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.02" eventid="1123" heatid="40046" lane="8">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:30.20" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.99" eventid="1163" heatid="40117" lane="7">
                  <MEETINFO name="DMS 2. Landesliga SHSV" city="Kiel" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:02:52.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.66" eventid="1207" heatid="40162" lane="2">
                  <MEETINFO name="SHSV-Sprintmehrkampf &amp; Staffel-MS" city="Lübeck" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:42.66" />
                </ENTRY>
                <ENTRY entrytime="00:05:18.90" eventid="1247" heatid="40239" lane="4">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:05:07.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.02" eventid="1267" heatid="40279" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:04.42" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.84" eventid="1307" heatid="40355" lane="8">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:42.11" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.86" eventid="1347" heatid="40415" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:21.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.55" eventid="1387" heatid="40477" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:01:16.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4736" nation="GER" region="04" clubid="35375" name="PSV Cottbus 90">
          <ATHLETES>
            <ATHLETE firstname="Nils" lastname="Wank" birthdate="2014-01-01" gender="M" nation="GER" license="448458" athleteid="35556">
              <ENTRIES>
                <ENTRY entrytime="00:11:15.00" eventid="1093" heatid="40013" lane="7" />
                <ENTRY entrytime="00:00:33.23" eventid="1133" heatid="40066" lane="2">
                  <MEETINFO name="16. Internationales Nachwuchsschwimmfest" city="Cottbus" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:33.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.93" eventid="1173" heatid="40132" lane="7">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:02:58.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.25" eventid="1217" heatid="40176" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:44.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.98" eventid="1237" heatid="40220" lane="4">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:19.12" />
                </ENTRY>
                <ENTRY entrytime="00:05:33.70" eventid="1257" heatid="40249" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:05:26.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.79" eventid="1277" heatid="40292" lane="3">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:12.27" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.29" eventid="1317" heatid="40365" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:55.41" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.85" eventid="1357" heatid="40424" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:32.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.34" eventid="1397" heatid="40487" lane="1">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:01:37.34" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fabian" lastname="Scherret" birthdate="2014-01-01" gender="M" nation="GER" license="448455" athleteid="35523">
              <ENTRIES>
                <ENTRY entrytime="00:11:15.00" eventid="1093" heatid="40013" lane="2" />
                <ENTRY entrytime="00:00:34.59" eventid="1133" heatid="40063" lane="5">
                  <MEETINFO name="16. Internationales Nachwuchsschwimmfest" city="Cottbus" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:34.59" />
                </ENTRY>
                <ENTRY entrytime="00:03:26.77" eventid="1153" heatid="40103" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:03:15.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.96" eventid="1217" heatid="40178" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:42.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.86" eventid="1237" heatid="40217" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:22.97" />
                </ENTRY>
                <ENTRY entrytime="00:05:52.43" eventid="1257" heatid="40247" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:05:52.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.33" eventid="1277" heatid="40290" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:16.81" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.50" eventid="1317" heatid="40364" lane="3">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:03:04.56" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.33" eventid="1357" heatid="40422" lane="6">
                  <MEETINFO name="Piranha Meeting" city="Hannover" course="LCM" approved="GER" date="2025-03-01" qualificationtime="00:02:56.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.89" eventid="1377" heatid="40461" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:39.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Niklas" lastname="Thierfelder" birthdate="2011-01-01" gender="M" nation="GER" license="424705" athleteid="35534">
              <ENTRIES>
                <ENTRY entrytime="00:05:35.00" eventid="1073" heatid="40000" lane="2" />
                <ENTRY entrytime="00:19:45.00" eventid="1113" heatid="40024" lane="6" />
                <ENTRY entrytime="00:02:55.26" eventid="1153" heatid="40107" lane="3">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:45.10" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.24" eventid="1173" heatid="40140" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:16.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.65" eventid="1197" heatid="40153" lane="5">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:02:29.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.05" eventid="1237" heatid="40230" lane="6">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:04.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.43" eventid="1277" heatid="40304" lane="4">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:01:00.43" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.58" eventid="1317" heatid="40373" lane="2">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:02:27.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.17" eventid="1377" heatid="40472" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:28.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.77" eventid="1397" heatid="40493" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:03.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Thomas" birthdate="2014-01-01" gender="M" nation="GER" license="448478" athleteid="35545">
              <ENTRIES>
                <ENTRY entrytime="00:06:20.00" eventid="1073" heatid="39998" lane="2" />
                <ENTRY entrytime="00:22:00.00" eventid="1113" heatid="40022" lane="3" />
                <ENTRY entrytime="00:00:31.82" eventid="1133" heatid="40069" lane="6">
                  <MEETINFO name="Talentewettkampf" city="Cottbus" course="SCM" approved="GER" date="2025-06-22" qualificationtime="00:00:31.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.66" eventid="1173" heatid="40134" lane="5">
                  <MEETINFO name="Piranha Meeting" city="Hannover" course="LCM" approved="GER" date="2025-03-02" qualificationtime="00:02:49.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.17" eventid="1197" heatid="40152" lane="2">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:02:56.17" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.49" eventid="1257" heatid="40252" lane="3">
                  <MEETINFO name="Norddeutsche Mehrkampfmeisterschaften" city="Bremen" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:05:15.49" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.96" eventid="1277" heatid="40296" lane="7">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:01:09.96" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.91" eventid="1317" heatid="40368" lane="2">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:02:46.78" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.88" eventid="1357" heatid="40426" lane="6">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:32.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.36" eventid="1397" heatid="40489" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:21.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nora" lastname="Kretzschmar" birthdate="2014-01-01" gender="F" nation="GER" license="448459" athleteid="35470">
              <ENTRIES>
                <ENTRY entrytime="00:22:15.00" eventid="1103" heatid="40020" lane="4" />
                <ENTRY entrytime="00:00:36.34" eventid="1123" heatid="40028" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:34.66" />
                </ENTRY>
                <ENTRY entrytime="00:03:35.08" eventid="1143" heatid="40090" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:03:17.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.34" eventid="1207" heatid="40158" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:43.94" />
                </ENTRY>
                <ENTRY entrytime="00:05:51.72" eventid="1247" heatid="40235" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:05:40.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.92" eventid="1267" heatid="40263" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:14.84" />
                </ENTRY>
                <ENTRY entrytime="00:03:14.53" eventid="1307" heatid="40349" lane="7">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:03:10.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.80" eventid="1327" heatid="40379" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:36.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.22" eventid="1347" heatid="40406" lane="2">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:46.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:46.00" eventid="1387" heatid="40475" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Joe" lastname="Betker" birthdate="2007-01-01" gender="M" nation="GER" license="366280" athleteid="35376">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.00" eventid="1133" heatid="40079" lane="6" />
                <ENTRY entrytime="00:00:36.00" eventid="1217" heatid="40184" lane="3" />
                <ENTRY entrytime="00:01:15.00" eventid="1237" heatid="40225" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="1277" heatid="40306" lane="1" />
                <ENTRY entrytime="00:00:32.00" eventid="1297" heatid="40339" lane="7" />
                <ENTRY entrytime="00:01:20.00" eventid="1337" heatid="40399" lane="1" />
                <ENTRY entrytime="00:00:34.00" eventid="1377" heatid="40469" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Til" lastname="Betker" birthdate="2010-01-01" gender="M" nation="GER" license="412412" athleteid="35384">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.11" eventid="1133" heatid="40082" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:26.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.31" eventid="1153" heatid="40108" lane="3">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:02:51.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.91" eventid="1217" heatid="40186" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:33.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.41" eventid="1237" heatid="40229" lane="8">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:01:10.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.01" eventid="1277" heatid="40304" lane="1">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:00.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.90" eventid="1297" heatid="40341" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:28.16" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.80" eventid="1337" heatid="40400" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:14.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.00" eventid="1377" heatid="40469" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:30.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.75" eventid="1397" heatid="40493" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:04.50" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Bastian" lastname="Welach" birthdate="2013-01-01" gender="M" nation="GER" license="444440" athleteid="35567">
              <ENTRIES>
                <ENTRY entrytime="00:06:10.00" eventid="1073" heatid="39998" lane="4" />
                <ENTRY entrytime="00:21:00.00" eventid="1113" heatid="40023" lane="3" />
                <ENTRY entrytime="00:00:31.35" eventid="1133" heatid="40070" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:30.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.86" eventid="1173" heatid="40134" lane="1">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:48.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.65" eventid="1237" heatid="40222" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:16.16" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.09" eventid="1257" heatid="40252" lane="5">
                  <MEETINFO name="Norddeutsche Mehrkampfmeisterschaften" city="Bremen" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:05:15.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.33" eventid="1277" heatid="40297" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:06.99" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.79" eventid="1317" heatid="40366" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:51.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.70" eventid="1357" heatid="40427" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:22.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.22" eventid="1377" heatid="40466" lane="2">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:35.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.02" eventid="1397" heatid="40489" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:15.22" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ida" lastname="Kretzschmar" birthdate="2011-01-01" gender="F" nation="GER" license="424712" athleteid="35464">
              <ENTRIES>
                <ENTRY entrytime="00:11:00.00" eventid="1083" heatid="40007" lane="5" />
                <ENTRY entrytime="00:00:30.91" eventid="1123" heatid="40046" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:30.27" />
                </ENTRY>
                <ENTRY entrytime="00:03:04.20" eventid="1143" heatid="40096" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:56.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.27" eventid="1207" heatid="40169" lane="5">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:36.86" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.00" eventid="1247" heatid="40240" lane="4" />
                <ENTRY entrytime="00:01:09.08" eventid="1267" heatid="40275" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:05.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.68" eventid="1327" heatid="40387" lane="2">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:20.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.60" eventid="1347" heatid="40415" lane="3">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:20.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.68" eventid="1367" heatid="40452" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:35.68" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lilly" lastname="Dommach" birthdate="2013-01-01" gender="F" nation="GER" license="444666" athleteid="35394">
              <ENTRIES>
                <ENTRY entrytime="00:06:09.76" eventid="1063" heatid="39994" lane="3" />
                <ENTRY entrytime="00:21:45.00" eventid="1103" heatid="40021" lane="8" />
                <ENTRY entrytime="00:00:31.49" eventid="1123" heatid="40043" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:30.63" />
                </ENTRY>
                <ENTRY entrytime="00:03:10.69" eventid="1143" heatid="40094" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:03:02.82" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.97" eventid="1187" heatid="40148" lane="3">
                  <MEETINFO name="Norddeutsche Mehrkampfmeisterschaften" city="Bremen" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:02:54.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.11" eventid="1207" heatid="40166" lane="2">
                  <MEETINFO name="Talentewettkampf" city="Cottbus" course="SCM" approved="GER" date="2025-06-22" qualificationtime="00:00:37.06" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.40" eventid="1247" heatid="40240" lane="3">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:15.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.06" eventid="1287" heatid="40323" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:32.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.25" eventid="1327" heatid="40385" lane="4">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:25.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.18" eventid="1347" heatid="40413" lane="1">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:28.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.81" eventid="1387" heatid="40481" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:15.97" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Frieda" lastname="Medwesch" birthdate="2014-01-01" gender="F" nation="GER" license="448461" athleteid="35487">
              <ENTRIES>
                <ENTRY entrytime="00:06:20.00" eventid="1063" heatid="39994" lane="1" />
                <ENTRY entrytime="00:22:15.00" eventid="1103" heatid="40020" lane="5" />
                <ENTRY entrytime="00:00:32.31" eventid="1123" heatid="40038" lane="8">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:31.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:57.48" eventid="1163" heatid="40117" lane="1">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:54.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.12" eventid="1227" heatid="40198" lane="3">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:21.23" />
                </ENTRY>
                <ENTRY entrytime="00:05:22.36" eventid="1247" heatid="40238" lane="4">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:05:20.39" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.11" eventid="1267" heatid="40271" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:09.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.26" eventid="1287" heatid="40316" lane="1">
                  <MEETINFO name="Talentewettkampf" city="Cottbus" course="SCM" approved="GER" date="2025-06-22" qualificationtime="00:00:36.11" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.41" eventid="1307" heatid="40355" lane="1">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-08" qualificationtime="00:02:52.41" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.50" eventid="1347" heatid="40412" lane="6">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:31.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.22" eventid="1387" heatid="40478" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:22.55" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anton" lastname="Freitag" birthdate="2014-01-01" gender="M" nation="GER" license="448481" athleteid="35406">
              <ENTRIES>
                <ENTRY entrytime="00:06:20.00" eventid="1073" heatid="39998" lane="6" />
                <ENTRY entrytime="00:11:15.00" eventid="1093" heatid="40013" lane="6" />
                <ENTRY entrytime="00:00:35.13" eventid="1133" heatid="40063" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:33.80" />
                </ENTRY>
                <ENTRY entrytime="00:03:15.89" eventid="1173" heatid="40129" lane="6">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:03:15.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.99" eventid="1217" heatid="40175" lane="8">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:48.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.00" eventid="1237" heatid="40215" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:28.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.29" eventid="1277" heatid="40289" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:14.46" />
                </ENTRY>
                <ENTRY entrytime="00:03:19.35" eventid="1317" heatid="40362" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:03:06.11" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.52" eventid="1357" heatid="40422" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:39.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:47.00" eventid="1397" heatid="40486" lane="2">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:01:50.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fritz" lastname="Kaiser" birthdate="2014-01-01" gender="M" nation="GER" license="448472" athleteid="35441">
              <ENTRIES>
                <ENTRY entrytime="00:06:20.00" eventid="1073" heatid="39998" lane="5" />
                <ENTRY entrytime="00:21:12.13" eventid="1113" heatid="40023" lane="7">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:21:12.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.94" eventid="1133" heatid="40067" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:32.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.88" eventid="1173" heatid="40132" lane="2">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:49.02" />
                </ENTRY>
                <ENTRY entrytime="00:03:11.40" eventid="1197" heatid="40151" lane="4">
                  <MEETINFO name="Piranha Meeting" city="Hannover" course="LCM" approved="GER" date="2025-03-01" qualificationtime="00:03:11.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.39" eventid="1237" heatid="40219" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:22.81" />
                </ENTRY>
                <ENTRY entrytime="00:05:20.57" eventid="1257" heatid="40251" lane="6">
                  <MEETINFO name="Norddeutsche Mehrkampfmeisterschaften" city="Bremen" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:05:20.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.03" eventid="1297" heatid="40333" lane="1">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:36.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.47" eventid="1317" heatid="40366" lane="4">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:52.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.46" eventid="1357" heatid="40426" lane="4">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:32.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.73" eventid="1397" heatid="40488" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:21.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Estella" lastname="Greif" birthdate="2013-01-01" gender="F" nation="GER" license="444439" athleteid="35417">
              <ENTRIES>
                <ENTRY entrytime="00:06:05.54" eventid="1063" heatid="39995" lane="8" />
                <ENTRY entrytime="00:21:28.08" eventid="1103" heatid="40021" lane="7" />
                <ENTRY entrytime="00:00:30.17" eventid="1123" heatid="40049" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:28.34" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.97" eventid="1143" heatid="40097" lane="1">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:03:01.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.43" eventid="1207" heatid="40167" lane="5">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:36.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.48" eventid="1227" heatid="40208" lane="8">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:09.11" />
                </ENTRY>
                <ENTRY entrytime="00:04:58.87" eventid="1247" heatid="40243" lane="2">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:04:58.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.71" eventid="1267" heatid="40278" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:03.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.17" eventid="1307" heatid="40357" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:37.80" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.76" eventid="1347" heatid="40415" lane="6">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:20.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.02" eventid="1387" heatid="40478" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:18.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Sachs" birthdate="2013-01-01" gender="M" nation="GER" license="444445" athleteid="35499">
              <ENTRIES>
                <ENTRY entrytime="00:06:10.00" eventid="1073" heatid="39999" lane="1" />
                <ENTRY entrytime="00:21:00.00" eventid="1113" heatid="40023" lane="6" />
                <ENTRY entrytime="00:00:30.90" eventid="1133" heatid="40071" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:28.99" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.58" eventid="1173" heatid="40137" lane="1">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:02:40.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.69" eventid="1237" heatid="40226" lane="5">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:01:13.69" />
                </ENTRY>
                <ENTRY entrytime="00:05:18.02" eventid="1257" heatid="40252" lane="8">
                  <MEETINFO name="Norddeutsche Mehrkampfmeisterschaften" city="Bremen" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:05:18.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.21" eventid="1277" heatid="40296" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:05.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.05" eventid="1317" heatid="40369" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:40.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.60" eventid="1357" heatid="40427" lane="8">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:26.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.35" eventid="1397" heatid="40489" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:14.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Finn" lastname="Jentsch" birthdate="2014-01-01" gender="M" nation="GER" license="448470" athleteid="35429">
              <ENTRIES>
                <ENTRY entrytime="00:06:20.00" eventid="1073" heatid="39998" lane="3" />
                <ENTRY entrytime="00:22:00.00" eventid="1113" heatid="40022" lane="5" />
                <ENTRY entrytime="00:00:32.98" eventid="1133" heatid="40067" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:31.86" />
                </ENTRY>
                <ENTRY entrytime="00:03:16.43" eventid="1153" heatid="40104" lane="7">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:03:10.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.83" eventid="1217" heatid="40177" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:41.47" />
                </ENTRY>
                <ENTRY entrytime="00:05:36.34" eventid="1257" heatid="40248" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:05:17.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.66" eventid="1277" heatid="40293" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:12.29" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.86" eventid="1317" heatid="40364" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:50.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.10" eventid="1337" heatid="40394" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:31.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.53" eventid="1357" heatid="40424" lane="3">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:36.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.96" eventid="1397" heatid="40486" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lina-Luisa" lastname="Sagroda" birthdate="2014-01-01" gender="F" nation="GER" license="448475" athleteid="35510">
              <ENTRIES>
                <ENTRY entrytime="00:06:20.00" eventid="1063" heatid="39994" lane="7" />
                <ENTRY entrytime="00:22:15.00" eventid="1103" heatid="40020" lane="3" />
                <ENTRY entrytime="00:00:33.56" eventid="1123" heatid="40033" lane="4">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:32.63" />
                </ENTRY>
                <ENTRY entrytime="00:03:19.32" eventid="1143" heatid="40093" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:03:07.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.37" eventid="1207" heatid="40164" lane="7">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:39.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.41" eventid="1227" heatid="40197" lane="2">
                  <MEETINFO name="16. Internationales Nachwuchsschwimmfest" city="Cottbus" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:25.41" />
                </ENTRY>
                <ENTRY entrytime="00:05:37.87" eventid="1247" heatid="40237" lane="8">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:05:37.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.05" eventid="1267" heatid="40267" lane="8">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:14.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:57.79" eventid="1307" heatid="40352" lane="5">
                  <MEETINFO name="Winterschwimmfest" city="Cottbus" course="SCM" approved="GER" date="2025-02-22" qualificationtime="00:02:57.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.57" eventid="1327" heatid="40383" lane="5">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:27.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.30" eventid="1347" heatid="40410" lane="8">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:36.11" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.31" eventid="1387" heatid="40476" lane="2">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:26.74" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Liebig" birthdate="2013-01-01" gender="M" nation="GER" license="444456" athleteid="35476">
              <ENTRIES>
                <ENTRY entrytime="00:06:10.00" eventid="1073" heatid="39999" lane="8" />
                <ENTRY entrytime="00:21:00.00" eventid="1113" heatid="40023" lane="2" />
                <ENTRY entrytime="00:00:33.09" eventid="1133" heatid="40066" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:31.80" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.90" eventid="1173" heatid="40133" lane="1">
                  <MEETINFO name="16. Internationales Nachwuchsschwimmfest" city="Cottbus" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:54.90" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.15" eventid="1237" heatid="40221" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:15.53" />
                </ENTRY>
                <ENTRY entrytime="00:05:19.13" eventid="1257" heatid="40251" lane="5">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:05:19.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.44" eventid="1277" heatid="40294" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:09.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.64" eventid="1317" heatid="40367" lane="2">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:02:42.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.59" eventid="1357" heatid="40427" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:28.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.18" eventid="1397" heatid="40489" lane="5">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:16.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Martins" lastname="Zabothens" birthdate="2005-01-01" gender="M" nation="GER" license="342627" athleteid="36376">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.50" eventid="1297" heatid="40347" lane="1">
                  <MEETINFO name="Sprintertag" city="Chemnitz" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:25.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.50" eventid="1397" heatid="40496" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Benjamin Robin" lastname="Klausch" birthdate="2010-01-01" gender="M" nation="GER" license="412416" athleteid="35453">
              <ENTRIES>
                <ENTRY entrytime="00:05:23.83" eventid="1073" heatid="40000" lane="6" />
                <ENTRY entrytime="00:19:15.00" eventid="1113" heatid="40024" lane="4" />
                <ENTRY entrytime="00:00:25.85" eventid="1133" heatid="40086" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:25.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.50" eventid="1173" heatid="40140" lane="8">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:02:19.61" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.01" eventid="1217" heatid="40184" lane="2">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:00:36.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.26" eventid="1237" heatid="40230" lane="5">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:03.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.87" eventid="1277" heatid="40308" lane="4">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:00:56.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.04" eventid="1337" heatid="40399" lane="8">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:01:20.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.69" eventid="1377" heatid="40473" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:28.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.02" eventid="1397" heatid="40494" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:03.08" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.37" eventid="1185" heatid="40146" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="35534" number="1" />
                    <RELAYPOSITION athleteid="35384" number="2" />
                    <RELAYPOSITION athleteid="35453" number="3" />
                    <RELAYPOSITION athleteid="35376" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <ENTRIES>
                <ENTRY entrytime="00:02:24.40" eventid="1185" heatid="40145" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="35499" number="1" />
                    <RELAYPOSITION athleteid="35429" number="2" />
                    <RELAYPOSITION athleteid="35545" number="3" />
                    <RELAYPOSITION athleteid="35567" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <ENTRIES>
                <ENTRY entrytime="00:02:13.26" eventid="1183" heatid="40144" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="35417" number="1" />
                    <RELAYPOSITION athleteid="35464" number="2" />
                    <RELAYPOSITION athleteid="35394" number="3" />
                    <RELAYPOSITION athleteid="35487" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="3513" nation="GER" region="14" clubid="34877" name="SV Wiking Kiel">
          <ATHLETES>
            <ATHLETE firstname="Alexander" lastname="Wieland" birthdate="2014-01-01" gender="M" nation="GER" license="462629" athleteid="34922">
              <ENTRIES>
                <ENTRY entrytime="00:11:14.00" eventid="1093" heatid="40013" lane="5">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:11:54.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.24" eventid="1133" heatid="40064" lane="6">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:33.28" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.10" eventid="1173" heatid="40131" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:03:01.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.56" eventid="1237" heatid="40219" lane="5">
                  <MEETINFO name="31. Herbst-Nachwuchsmeeting" city="Kiel" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:01:24.56" />
                </ENTRY>
                <ENTRY entrytime="00:05:51.99" eventid="1257" heatid="40247" lane="4">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:05:51.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.96" eventid="1297" heatid="40334" lane="2">
                  <MEETINFO name="SHSV-Sprintmehrkampf &amp; Staffel-MS" city="Lübeck" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:35.96" />
                </ENTRY>
                <ENTRY entrytime="00:03:09.49" eventid="1317" heatid="40364" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:03:09.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.86" eventid="1377" heatid="40463" lane="2">
                  <MEETINFO name="31. Herbst-Nachwuchsmeeting" city="Kiel" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:39.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.41" eventid="1397" heatid="40488" lane="1">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:28.22" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jolie" lastname="Sobottka" birthdate="2008-01-01" gender="F" nation="GER" license="404150" athleteid="34907">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.06" eventid="1123" heatid="40056" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:28.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.34" eventid="1163" heatid="40125" lane="5">
                  <MEETINFO name="DMS 2. Landesliga SHSV" city="Kiel" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:02:35.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.19" eventid="1227" heatid="40212" lane="7">
                  <MEETINFO name="32. Sommerwettkämpfe mit dem 1. Kieler-Woche-Pokal" city="Kiel" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:10.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.62" eventid="1267" heatid="40285" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:01.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.47" eventid="1287" heatid="40322" lane="7">
                  <MEETINFO name="1. Swim-Cup powered by Stadtwerke Solingen" city="Solingen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:33.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.10" eventid="1367" heatid="40458" lane="5">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:32.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Simon" lastname="Ludewigsen" birthdate="2011-01-01" gender="M" nation="GER" license="424986" athleteid="34886">
              <ENTRIES>
                <ENTRY entrytime="00:05:35.00" eventid="1073" heatid="40000" lane="7">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:05:35.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.56" eventid="1133" heatid="40074" lane="5">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:28.68" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.15" eventid="1153" heatid="40108" lane="4">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:49.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.47" eventid="1217" heatid="40185" lane="2">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:35.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.81" eventid="1237" heatid="40226" lane="3">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:13.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.00" eventid="1277" heatid="40299" lane="5">
                  <MEETINFO name="32. Sommerwettkämpfe mit dem 1. Kieler-Woche-Pokal" city="Kiel" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:05.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.54" eventid="1317" heatid="40371" lane="3">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:36.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.46" eventid="1337" heatid="40401" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:16.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.48" eventid="1377" heatid="40467" lane="6">
                  <MEETINFO name="SHSV-MS, JG-MS und SMK" city="Kiel" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:00:35.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.59" eventid="1397" heatid="40491" lane="5">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:10.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Sturm" birthdate="2012-01-01" gender="M" nation="GER" license="446482" athleteid="34914">
              <ENTRIES>
                <ENTRY entrytime="00:10:25.34" eventid="1093" heatid="40016" lane="7">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:10:11.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.11" eventid="1153" heatid="40108" lane="2">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:45.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.77" eventid="1217" heatid="40185" lane="8">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:35.77" />
                </ENTRY>
                <ENTRY entrytime="00:04:50.47" eventid="1257" heatid="40255" lane="4">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:04:50.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.44" eventid="1277" heatid="40300" lane="2">
                  <MEETINFO name="32. Sommerwettkämpfe mit dem 1. Kieler-Woche-Pokal" city="Kiel" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:04.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.86" eventid="1337" heatid="40400" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:17.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.92" eventid="1357" heatid="40431" lane="7">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:18.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Ludewigsen" birthdate="2013-01-01" gender="M" nation="GER" license="428696" athleteid="34878">
              <ENTRIES>
                <ENTRY entrytime="00:10:24.00" eventid="1093" heatid="40016" lane="2">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:11:38.45" />
                </ENTRY>
                <ENTRY entrytime="00:03:17.27" eventid="1153" heatid="40104" lane="1">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:03:12.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.68" eventid="1237" heatid="40220" lane="6">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:21.16" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.89" eventid="1277" heatid="40292" lane="6">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:01:12.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.85" eventid="1317" heatid="40365" lane="6">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:58.21" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.99" eventid="1337" heatid="40394" lane="4">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:31.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.92" eventid="1377" heatid="40464" lane="3">
                  <MEETINFO name="32. Sommerwettkämpfe mit dem 1. Kieler-Woche-Pokal" city="Kiel" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:37.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nele" lastname="Petersen" birthdate="2010-01-01" gender="F" nation="GER" license="421793" athleteid="34897">
              <ENTRIES>
                <ENTRY entrytime="00:10:44.00" eventid="1083" status="WDR" heatid="40009" lane="1" />
                <ENTRY entrytime="00:00:31.11" eventid="1123" heatid="40045" lane="8">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:30.81" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.00" eventid="1163" heatid="40119" lane="4">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:57.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.51" eventid="1227" heatid="40202" lane="5">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:20.51" />
                </ENTRY>
                <ENTRY entrytime="00:05:00.00" eventid="1247" heatid="40243" lane="1" />
                <ENTRY entrytime="00:01:08.19" eventid="1267" heatid="40277" lane="2">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:08.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.00" eventid="1287" heatid="40316" lane="3">
                  <MEETINFO name="32. Wiking-Pokal" city="Kiel" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:37.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.45" eventid="1347" heatid="40412" lane="3">
                  <MEETINFO name="50. Internationaler Förde - Pokal" city="Flensburg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:02:33.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.40" eventid="1367" heatid="40448" lane="6">
                  <MEETINFO name="Kreismeisterschaften" city="Kiel" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:36.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LVIV" nation="UKR" clubid="36720" name="LVIV Sports School of Sydoruk">
          <CONTACT email="rivak.kristi@gmail.com, sportschool.sydoruka@gmail" name="LVIV Sports School of Sydoruk" phone="+38 (096) 725-74-28" street="10 V.Yaneva Street, Lviv" zip="79000" />
          <ATHLETES>
            <ATHLETE firstname="Dmytro" lastname="Markiv" birthdate="2015-10-29" gender="M" nation="UKR" athleteid="36797">
              <ENTRIES>
                <ENTRY entrytime="00:03:42.98" entrycourse="LCM" eventid="1153" heatid="40102" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:00:46.49" entrycourse="LCM" eventid="1217" heatid="40175" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:43.49" entrycourse="LCM" eventid="1297" heatid="40331" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:01:45.99" entrycourse="LCM" eventid="1337" heatid="40391" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:03:03.99" entrycourse="LCM" eventid="1357" heatid="40421" lane="4">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Solomiia" lastname="Lytvyn" birthdate="2010-05-27" gender="F" nation="UKR" athleteid="36733">
              <ENTRIES>
                <ENTRY entrytime="00:10:44.20" entrycourse="LCM" eventid="1083" heatid="40009" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:00:31.80" entrycourse="LCM" eventid="1123" heatid="40041" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:01:18.30" entrycourse="LCM" eventid="1227" heatid="40205" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:01:09.67" entrycourse="LCM" eventid="1267" heatid="40273" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:02:49.80" entrycourse="LCM" eventid="1307" heatid="40356" lane="7">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lev" lastname="Dratver" birthdate="2015-07-22" gender="M" nation="UKR" athleteid="36721">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.92" entrycourse="LCM" eventid="1133" heatid="40060" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:01:43.32" entrycourse="LCM" eventid="1237" heatid="40214" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:26.98" entrycourse="LCM" eventid="1277" heatid="40287" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:03:11.42" entrycourse="LCM" eventid="1357" heatid="40421" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:00:46.21" entrycourse="LCM" eventid="1377" heatid="40460" lane="4">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mariia" lastname="Puchak" birthdate="2012-08-24" gender="F" nation="UKR" athleteid="36821">
              <ENTRIES>
                <ENTRY entrytime="00:05:53.70" entrycourse="LCM" eventid="1247" heatid="40235" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:01:14.70" entrycourse="LCM" eventid="1267" heatid="40267" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:03:02.70" entrycourse="LCM" eventid="1307" heatid="40351" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:02:41.70" entrycourse="LCM" eventid="1347" heatid="40409" lane="1">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ihor" lastname="Petryna" birthdate="2009-02-06" gender="M" nation="UKR" athleteid="36803">
              <ENTRIES>
                <ENTRY entrytime="00:09:30.70" entrycourse="LCM" eventid="1093" heatid="40018" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:00:27.70" entrycourse="LCM" eventid="1133" heatid="40080" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:04:34.70" entrycourse="LCM" eventid="1257" heatid="40258" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:24.70" entrycourse="LCM" eventid="1317" heatid="40373" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:02:07.70" entrycourse="LCM" eventid="1357" heatid="40436" lane="6">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Danylo" lastname="Fylypiv" birthdate="2008-09-21" gender="M" nation="UKR" athleteid="36774">
              <ENTRIES>
                <ENTRY entrytime="00:08:41.00" entrycourse="LCM" eventid="1093" heatid="40019" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:04:07.00" entrycourse="LCM" eventid="1257" heatid="40260" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:26.85" entrycourse="LCM" eventid="1297" heatid="40346" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:01:58.00" entrycourse="LCM" eventid="1357" heatid="40438" lane="5">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Volodymyr" lastname="Pasichnyk" birthdate="2009-04-25" gender="M" nation="UKR" athleteid="36739">
              <ENTRIES>
                <ENTRY entrytime="00:02:21.00" entrycourse="LCM" eventid="1173" heatid="40141" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:01:03.00" entrycourse="LCM" eventid="1237" heatid="40231" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:00:28.00" entrycourse="LCM" eventid="1297" heatid="40344" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:00:28.00" entrycourse="LCM" eventid="1377" heatid="40474" lane="1">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Stefaniia" lastname="Hladkova" birthdate="2013-04-28" gender="F" nation="UKR" athleteid="36785">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.30" eventid="1123" heatid="40034" lane="3" />
                <ENTRY entrytime="00:00:45.00" eventid="1207" heatid="40159" lane="2" />
                <ENTRY entrytime="00:05:50.00" eventid="1247" heatid="40235" lane="5" />
                <ENTRY entrytime="00:00:34.00" eventid="1287" heatid="40320" lane="4" />
                <ENTRY entrytime="00:01:30.00" eventid="1387" heatid="40477" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Rostyslav" lastname="Romaniv" birthdate="2014-10-02" gender="M" nation="UKR" athleteid="36744">
              <ENTRIES>
                <ENTRY entrytime="00:10:36.70" entrycourse="LCM" eventid="1093" heatid="40015" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:05:27.70" entrycourse="LCM" eventid="1257" heatid="40250" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:03:05.00" entrycourse="LCM" eventid="1317" heatid="40364" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:01:25.70" entrycourse="LCM" eventid="1397" heatid="40488" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:03:37.00" eventid="1153" heatid="40102" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Olha" lastname="Kuzyk" birthdate="2011-11-13" gender="F" nation="UKR" athleteid="36791">
              <ENTRIES>
                <ENTRY entrytime="00:10:40.43" entrycourse="LCM" eventid="1083" heatid="40009" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:02:40.36" entrycourse="LCM" eventid="1163" heatid="40123" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:01:14.25" entrycourse="LCM" eventid="1227" heatid="40209" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:02:38.32" entrycourse="LCM" eventid="1307" heatid="40359" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:00:34.20" entrycourse="LCM" eventid="1367" heatid="40455" lane="7">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Yaroslav" lastname="Kopetchak" birthdate="2012-06-29" gender="M" nation="UKR" athleteid="36727">
              <ENTRIES>
                <ENTRY entrytime="00:09:50.70" entrycourse="LCM" eventid="1093" status="WDR" heatid="40017" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:02:44.70" entrycourse="LCM" eventid="1153" status="WDR" heatid="40109" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:04:53.70" entrycourse="LCM" eventid="1257" status="WDR" heatid="40255" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:02:29.70" entrycourse="LCM" eventid="1317" status="WDR">
                </ENTRY>
                <ENTRY entrytime="00:01:11.70" entrycourse="LCM" eventid="1397" status="WDR">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ruslan" lastname="Rodevych" birthdate="2014-05-08" gender="M" nation="UKR" athleteid="36826">
              <ENTRIES>
                <ENTRY entrytime="00:10:03.47" entrycourse="LCM" eventid="1093" heatid="40016" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:02:59.00" entrycourse="LCM" eventid="1173" heatid="40132" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:05:27.00" entrycourse="LCM" eventid="1257" heatid="40250" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:35.00" entrycourse="LCM" eventid="1297" heatid="40335" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:02:55.50" entrycourse="LCM" eventid="1317" heatid="40366" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:19.50" entrycourse="LCM" eventid="1397" heatid="40489" lane="6">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Yurii" lastname="Shlyakhetko" birthdate="2013-12-27" gender="M" nation="UKR" athleteid="36755">
              <ENTRIES>
                <ENTRY entrytime="00:11:14.01" entrycourse="LCM" eventid="1093" heatid="40013" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:32.52" entrycourse="LCM" eventid="1133" heatid="40068" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:02:53.67" entrycourse="LCM" eventid="1173" heatid="40133" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:05:23.59" entrycourse="LCM" eventid="1257" heatid="40250" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:01:11.03" entrycourse="LCM" eventid="1277" heatid="40295" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:02:31.49" entrycourse="LCM" eventid="1357" heatid="40427" lane="5">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Yeva-Mariia" lastname="Smachylo" birthdate="2011-10-14" gender="F" nation="UKR" athleteid="36762">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.70" entrycourse="LCM" eventid="1123" heatid="40036" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:05:33.70" entrycourse="SCM" eventid="1247" heatid="40237" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:01:12.70" entrycourse="LCM" eventid="1267" heatid="40269" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:37.70" entrycourse="LCM" eventid="1347" heatid="40410" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:00:36.70" entrycourse="LCM" eventid="1367" heatid="40449" lane="5">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Oleksandr" lastname="Runts" birthdate="2013-04-10" gender="M" nation="UKR" athleteid="36750">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.70" entrycourse="LCM" eventid="1133" heatid="40065" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:10.70" entrycourse="LCM" eventid="1277" heatid="40295" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:00:35.50" entrycourse="LCM" eventid="1297" heatid="40334" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:00:39.70" entrycourse="LCM" eventid="1377" heatid="40463" lane="5">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Dmytro" lastname="Fylypiv" birthdate="2011-10-02" gender="M" nation="UKR" athleteid="36779">
              <ENTRIES>
                <ENTRY entrytime="00:04:59.34" entrycourse="LCM" eventid="1073" heatid="40001" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:02:33.71" entrycourse="LCM" eventid="1153" heatid="40111" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:02:23.86" entrycourse="LCM" eventid="1197" heatid="40155" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:02:23.01" entrycourse="LCM" eventid="1317" heatid="40374" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:02:12.12" entrycourse="LCM" eventid="1357" heatid="40434" lane="6">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Armen" lastname="Parsadanian" birthdate="2011-07-30" gender="M" nation="UKR" athleteid="36809">
              <ENTRIES>
                <ENTRY entrytime="00:19:15.40" entrycourse="LCM" eventid="1113" heatid="40024" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:00:29.50" entrycourse="LCM" eventid="1133" status="WDR" heatid="40075" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:04:52.60" entrycourse="LCM" eventid="1257" heatid="40255" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:35.80" entrycourse="LCM" eventid="1317" heatid="40372" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:02:19.10" entrycourse="LCM" eventid="1357" heatid="40431" lane="1">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karen" lastname="Parsadanian" birthdate="2011-07-30" gender="M" nation="UKR" athleteid="36815">
              <ENTRIES>
                <ENTRY entrytime="00:09:50.01" entrycourse="LCM" eventid="1093" status="WDR" heatid="40017" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:02:30.00" entrycourse="LCM" eventid="1173" heatid="40139" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:01:11.00" entrycourse="LCM" eventid="1237" heatid="40228" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:04.40" entrycourse="LCM" eventid="1277" heatid="40300" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:02:15.20" entrycourse="LCM" eventid="1357" heatid="40432" lane="4">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maksym" lastname="Susol" birthdate="2012-03-14" gender="M" nation="UKR" athleteid="36768">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.30" entrycourse="LCM" eventid="1133" heatid="40078" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:01:14.70" entrycourse="LCM" eventid="1237" heatid="40226" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:01:06.70" entrycourse="LCM" eventid="1277" heatid="40298" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:34.00" entrycourse="LCM" eventid="1337" heatid="40394" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:02:18.70" entrycourse="LCM" eventid="1357" heatid="40431" lane="6">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5149" nation="GER" region="12" clubid="37860" name="SV 1919 Grimma">
          <ATHLETES>
            <ATHLETE firstname="Alessandro" lastname="Munari" birthdate="2013-01-01" gender="M" nation="GER" license="445022" athleteid="37861">
              <ENTRIES>
                <ENTRY entrytime="00:11:07.82" eventid="1093" heatid="40014" lane="8">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:11:07.82" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.82" eventid="1133" heatid="40069" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:31.82" />
                </ENTRY>
                <ENTRY entrytime="00:03:20.00" eventid="1153" heatid="40103" lane="5" />
                <ENTRY entrytime="00:00:44.39" eventid="1217" heatid="40177" lane="2">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:44.39" />
                </ENTRY>
                <ENTRY entrytime="00:05:12.63" eventid="1257" heatid="40252" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:05:12.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.15" eventid="1317" heatid="40367" lane="8">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:55.15" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.08" eventid="1337" heatid="40394" lane="8">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:01:35.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.61" eventid="1357" heatid="40426" lane="7">
                  <MEETINFO name="29. Sparkassencup" city="Grimma" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:02:30.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.99" eventid="1397" heatid="40487" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:30.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karl" lastname="von Thun" birthdate="2005-01-01" gender="M" nation="GER" license="329642" athleteid="37871">
              <ENTRIES>
                <ENTRY entrytime="00:08:32.67" eventid="1093" heatid="40019" lane="5">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:08:32.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.23" eventid="1153" heatid="40110" lane="6" />
                <ENTRY entrytime="00:00:34.19" eventid="1217" heatid="40186" lane="6" />
                <ENTRY entrytime="00:01:02.68" eventid="1237" heatid="40231" lane="5">
                  <MEETINFO name="29. Sparkassencup" city="Grimma" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:57.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="USK" nation="CZE" clubid="36711" name="Univerzitní sportovní klub Praha">
          <CONTACT city="Prague" email="jan.rehor@plavecky.club" name="Michal Cervinka" />
          <ATHLETES>
            <ATHLETE firstname="Matyas" lastname="Bazant" birthdate="2010-05-12" gender="M" nation="CZE" athleteid="36712">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.85" entrycourse="SCM" eventid="1133" heatid="40084" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:02:23.26" entrycourse="SCM" eventid="1173" heatid="40140" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:37.66" entrycourse="LCM" eventid="1217" heatid="40182" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:04:28.72" entrycourse="SCM" eventid="1257" heatid="40259" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:00:58.46" entrycourse="SCM" eventid="1277" heatid="40308" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:02:39.55" entrycourse="LCM" eventid="1317" heatid="40371" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:02:07.40" entrycourse="SCM" eventid="1357" heatid="40436" lane="3">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3356" nation="GER" region="12" clubid="38894" name="SC Riesa">
          <ATHLETES>
            <ATHLETE firstname="Jonas" lastname="Schäfer" birthdate="2013-01-01" gender="M" nation="GER" license="449096" athleteid="38902">
              <ENTRIES>
                <ENTRY entrytime="00:20:29.07" eventid="1113" heatid="40024" lane="1">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:20:29.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.06" eventid="1133" heatid="40072" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:29.73" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.77" eventid="1197" heatid="40153" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:02:52.77" />
                </ENTRY>
                <ENTRY entrytime="00:05:03.14" eventid="1257" heatid="40254" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:04:59.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.91" eventid="1277" heatid="40298" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:06.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.38" eventid="1317" heatid="40370" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:43.38" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.72" eventid="1357" heatid="40430" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:21.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ole" lastname="Mühlmann" birthdate="2013-01-01" gender="M" nation="GER" license="446953" athleteid="38895">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.77" eventid="1133" heatid="40071" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:30.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.85" eventid="1217" heatid="40180" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:38.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.56" eventid="1237" heatid="40221" lane="2">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:01:21.56" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.91" eventid="1317" heatid="40369" lane="2">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:02:45.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.76" eventid="1337" heatid="40396" lane="7">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:28.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.75" eventid="1397" heatid="40490" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:16.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="7328" nation="GER" region="16" clubid="36382" name="Freibadverein Bad Blankenburg">
          <ATHLETES>
            <ATHLETE firstname="Ferdinand" lastname="Döring" birthdate="2006-01-01" gender="M" nation="GER" license="354729" athleteid="36383">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.75" eventid="1133" heatid="40086" lane="4">
                  <MEETINFO name="Saalfelder Feengrottenpokal" city="Saalfeld" course="SCM" approved="GER" date="2025-01-25" qualificationtime="00:00:25.50" />
                </ENTRY>
                <ENTRY entrytime="00:04:44.83" eventid="1257" heatid="40256" lane="6" />
                <ENTRY entrytime="00:00:27.08" eventid="1297" heatid="40346" lane="1">
                  <MEETINFO name="Plauener Herbst- Mehrkampf" city="Plauen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:27.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.17" eventid="1397" heatid="40495" lane="1">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:00.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Claudia" lastname="Rabold" birthdate="1975-01-01" gender="F" nation="GER" license="86089" athleteid="36388">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.04" eventid="1287" heatid="40318" lane="8">
                  <MEETINFO name="Saalfelder Feengrottenpokal" city="Saalfeld" course="SCM" approved="GER" date="2025-01-25" qualificationtime="00:00:35.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.29" eventid="1367" heatid="40453" lane="1">
                  <MEETINFO name="15. Deutsche Kurzbahnmeisterschaft der Masters" city="Essen" course="SCM" approved="GER" date="2025-11-29" qualificationtime="00:00:34.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lina" lastname="Reiher" birthdate="2006-01-01" gender="F" nation="GER" license="365728" athleteid="36396">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.95" eventid="1123" heatid="40040" lane="2">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:30.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.74" eventid="1227" heatid="40203" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:18.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.85" eventid="1267" heatid="40272" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:08.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.82" eventid="1367" heatid="40451" lane="6">
                  <MEETINFO name="Saalfelder Feengrottenpokal" city="Saalfeld" course="SCM" approved="GER" date="2025-01-25" qualificationtime="00:00:35.50" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Janik" lastname="Reiher" birthdate="2003-01-01" gender="M" nation="GER" license="298654" athleteid="36391">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.18" eventid="1133" heatid="40088" lane="4">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:23.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.78" eventid="1237" heatid="40231" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:59.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.30" eventid="1297" heatid="40345" lane="3">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:26.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.16" eventid="1377" heatid="40473" lane="6">
                  <MEETINFO name="15. Deutsche Kurzbahnmeisterschaft der Masters" city="Essen" course="SCM" approved="GER" date="2025-11-29" qualificationtime="00:00:27.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4344" nation="GER" region="02" clubid="34184" name="SV Augsburg 1911">
          <ATHLETES>
            <ATHLETE firstname="Leonie" lastname="von Bornstedt" birthdate="2014-01-01" gender="F" nation="GER" license="461018" athleteid="34804">
              <ENTRIES>
                <ENTRY entrytime="00:11:28.73" eventid="1083" heatid="40005" lane="6">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:11:49.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.66" eventid="1123" heatid="40026" lane="2" />
                <ENTRY entrytime="00:03:22.43" eventid="1143" heatid="40092" lane="6">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:03:20.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.74" eventid="1207" heatid="40162" lane="8">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:42.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.45" eventid="1227" heatid="40194" lane="7">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:26.15" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.26" eventid="1267" heatid="40266" lane="7">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:12.68" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.85" eventid="1327" heatid="40381" lane="3">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:29.60" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.53" eventid="1347" heatid="40407" lane="8">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:43.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.03" eventid="1367" heatid="40443" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Liana Emma" lastname="Koch" birthdate="2013-01-01" gender="F" nation="GER" license="448682" athleteid="34735">
              <ENTRIES>
                <ENTRY entrytime="00:05:53.19" eventid="1063" heatid="39995" lane="5">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:05:39.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.03" eventid="1123" heatid="40045" lane="4">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:30.48" />
                </ENTRY>
                <ENTRY entrytime="00:03:09.13" eventid="1163" heatid="40114" lane="1">
                  <MEETINFO name="Regionale Bestenkämpfe - Nord" city="Augsburg" course="SCM" approved="GER" date="2025-03-16" qualificationtime="00:02:50.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.30" eventid="1187" heatid="40149" lane="7">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:38.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.95" eventid="1227" heatid="40196" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:14.79" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.39" eventid="1267" heatid="40277" lane="1">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:06.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.12" eventid="1307" heatid="40356" lane="3">
                  <MEETINFO name="BaWü &amp; Süddt Meisterschaften SMK" city="Stuttgart" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:48.12" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.27" eventid="1347" heatid="40412" lane="4">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:30.68" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.14" eventid="1387" heatid="40482" lane="5">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:01:11.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Brummer" birthdate="2011-01-01" gender="F" nation="GER" license="423751" athleteid="34686">
              <ENTRIES>
                <ENTRY entrytime="00:10:03.06" eventid="1083" heatid="40010" lane="5">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:09:43.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.60" eventid="1123" heatid="40052" lane="1">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:00:29.60" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.45" eventid="1163" heatid="40125" lane="2">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:02:36.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.60" eventid="1187" heatid="40149" lane="3">
                  <MEETINFO name="Regionale Bestenkämpfe - Nord" city="Augsburg" course="SCM" approved="GER" date="2025-03-16" qualificationtime="00:02:42.10" />
                </ENTRY>
                <ENTRY entrytime="00:04:49.18" eventid="1247" heatid="40244" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:04:40.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.39" eventid="1267" heatid="40281" lane="5">
                  <MEETINFO name="Regionale Bestenkämpfe - Nord" city="Augsburg" course="SCM" approved="GER" date="2025-03-16" qualificationtime="00:01:02.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.76" eventid="1287" heatid="40326" lane="6">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:31.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.85" eventid="1347" heatid="40418" lane="1">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:16.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.34" eventid="1387" heatid="40484" lane="4">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:01:08.72" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Focke" birthdate="2014-01-01" gender="F" nation="GER" license="438386" athleteid="34706">
              <ENTRIES>
                <ENTRY entrytime="00:06:06.75" eventid="1063" heatid="39994" lane="4">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:05:50.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.57" eventid="1123" heatid="40031" lane="1" />
                <ENTRY entrytime="00:03:10.06" eventid="1143" heatid="40094" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:03:02.78" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.60" eventid="1187" heatid="40148" lane="6">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-11" qualificationtime="00:02:52.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.15" eventid="1227" heatid="40201" lane="2">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:18.20" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.26" eventid="1287" heatid="40320" lane="2">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:34.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.35" eventid="1327" heatid="40385" lane="6">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:24.17" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.11" eventid="1347" heatid="40411" lane="8">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:34.38" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.28" eventid="1387" heatid="40481" lane="2">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:01:16.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Vincent" lastname="Staudinger" birthdate="2012-01-01" gender="M" nation="GER" license="436775" athleteid="34784">
              <ENTRIES>
                <ENTRY entrytime="00:03:14.94" eventid="1153" heatid="40104" lane="3">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:03:00.14" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.72" eventid="1173" heatid="40137" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften" city="Bobingen" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:02:40.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.33" eventid="1237" heatid="40225" lane="8">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:13.67" />
                </ENTRY>
                <ENTRY entrytime="00:05:16.54" eventid="1257" heatid="40252" lane="7">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:05:12.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.33" eventid="1277" heatid="40298" lane="1">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:06.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.92" eventid="1337" heatid="40395" lane="4">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:24.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.29" eventid="1357" heatid="40428" lane="6">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:26.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.78" eventid="1377" heatid="40462" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Bögl" birthdate="2012-01-01" gender="F" nation="GER" license="441408" athleteid="34676">
              <ENTRIES>
                <ENTRY entrytime="00:10:48.27" eventid="1083" heatid="40008" lane="6">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:10:26.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.16" eventid="1123" heatid="40049" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:29.62" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.33" eventid="1143" heatid="40095" lane="6">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:03:00.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.94" eventid="1207" heatid="40170" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:36.64" />
                </ENTRY>
                <ENTRY entrytime="00:05:19.51" eventid="1247" heatid="40239" lane="6">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:05:06.69" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.02" eventid="1267" heatid="40279" lane="5">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:04.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.58" eventid="1287" heatid="40321" lane="4">
                  <MEETINFO name="Bezirksmeisterschaften" city="Bobingen" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:33.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.07" eventid="1347" heatid="40414" lane="4">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:20.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.57" eventid="1387" heatid="40480" lane="4">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:14.93" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Patrizia Yuexin" lastname="Stradovnik" birthdate="2011-01-01" gender="F" nation="BEL" license="478507" athleteid="34794">
              <ENTRIES>
                <ENTRY entrytime="00:18:45.61" eventid="1103" heatid="40021" lane="5">
                  <MEETINFO name="BaWü Meisterschaften (offene Klasse/Jugend A+B)" city="Freiburg" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:18:45.61" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.72" eventid="1123" heatid="40051" lane="2">
                  <MEETINFO name="BaWü Meisterschaften (offene Klasse/Jugend A+B)" city="Freiburg" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:00:29.72" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.83" eventid="1143" heatid="40096" lane="8">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-28" qualificationtime="00:03:05.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.11" eventid="1187" heatid="40150" lane="2">
                  <MEETINFO name="BaWü Meisterschaften (offene Klasse/Jugend A+B)" city="Freiburg" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:02:38.11" />
                </ENTRY>
                <ENTRY entrytime="00:04:47.30" eventid="1247" heatid="40244" lane="5">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:04:40.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.14" eventid="1267" heatid="40282" lane="2">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:01:04.14" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.74" eventid="1307" heatid="40359" lane="8">
                  <MEETINFO name="BaWü Meisterschaften (offene Klasse/Jugend A+B)" city="Freiburg" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:02:38.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.20" eventid="1347" heatid="40418" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:16.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.35" eventid="1387" heatid="40484" lane="8">
                  <MEETINFO name="International Sindelfingen Swimming Championship" city="Sindelfingen" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:01:11.35" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Nuber" birthdate="2015-01-01" gender="F" nation="GER" license="478573" athleteid="34774">
              <ENTRIES>
                <ENTRY entrytime="00:11:57.38" eventid="1083" heatid="40004" lane="1">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:12:12.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.53" eventid="1123" heatid="40026" lane="5">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:39.53" />
                </ENTRY>
                <ENTRY entrytime="00:03:11.24" eventid="1163" heatid="40113" lane="4">
                  <MEETINFO name="12. BSV Bezirksvergleich im Schwimmen" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:03:04.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.36" eventid="1227" heatid="40193" lane="7">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:31.75" />
                </ENTRY>
                <ENTRY entrytime="00:06:15.89" eventid="1247" heatid="40234" lane="6">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:06:15.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.83" eventid="1267" heatid="40261" lane="4">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:21.20" />
                </ENTRY>
                <ENTRY entrytime="00:03:11.60" eventid="1307" heatid="40349" lane="3">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-11" qualificationtime="00:03:11.60" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.50" eventid="1347" heatid="40405" lane="3">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:58.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.00" eventid="1387" heatid="40476" lane="3">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:35.76" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Kaminski" birthdate="2012-01-01" gender="F" nation="GER" license="448676" athleteid="34716">
              <ENTRIES>
                <ENTRY entrytime="00:10:48.32" eventid="1083" heatid="40008" lane="2">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:10:11.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.85" eventid="1123" heatid="40041" lane="6">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:30.79" />
                </ENTRY>
                <ENTRY entrytime="00:02:57.85" eventid="1143" heatid="40098" lane="1">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:02:52.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.15" eventid="1207" heatid="40168" lane="5">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:37.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.25" eventid="1227" heatid="40203" lane="7">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:15.37" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.79" eventid="1267" heatid="40273" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:07.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.00" eventid="1327" heatid="40388" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:21.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.86" eventid="1347" heatid="40415" lane="2">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:23.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.99" eventid="1367" heatid="40447" lane="6">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:37.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Elana" lastname="Moreira dos Santos" birthdate="2014-01-01" gender="F" nation="GER" license="449912" athleteid="34755">
              <ENTRIES>
                <ENTRY entrytime="00:11:03.97" eventid="1083" heatid="40006" lane="5">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:10:37.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.10" eventid="1123" heatid="40045" lane="7">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:00:31.10" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.91" eventid="1163" heatid="40118" lane="5">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:44.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.39" eventid="1227" heatid="40202" lane="8">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:01:17.15" />
                </ENTRY>
                <ENTRY entrytime="00:05:12.28" eventid="1247" heatid="40241" lane="5">
                  <MEETINFO name="BaWü &amp; Süddt Meisterschaften SMK" city="Stuttgart" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:05:12.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.13" eventid="1267" heatid="40275" lane="2">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:06.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.13" eventid="1307" heatid="40355" lane="3">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:47.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.95" eventid="1347" heatid="40415" lane="1">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:24.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.02" eventid="1387" heatid="40478" lane="2">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:21.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Srecko" lastname="Nikolic" birthdate="2009-01-01" gender="M" nation="GER" license="482303" athleteid="34765">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.18" eventid="1133" heatid="40079" lane="1">
                  <MEETINFO name="2. SUN-SWIM Trophy" city="Neckarsulm" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:00:28.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.05" eventid="1153" heatid="40108" lane="5">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:45.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.00" eventid="1217" heatid="40183" lane="1" />
                <ENTRY entrytime="00:01:14.23" eventid="1237" heatid="40226" lane="2">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:07.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.51" eventid="1277" heatid="40306" lane="5">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:59.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.99" eventid="1337" heatid="40400" lane="5">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:16.99" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.13" eventid="1357" heatid="40432" lane="1">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:16.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.59" eventid="1377" heatid="40467" lane="7" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Meyer" birthdate="2012-01-01" gender="M" nation="GER" license="442163" athleteid="34745">
              <ENTRIES>
                <ENTRY entrytime="00:10:19.98" eventid="1093" heatid="40016" lane="3" />
                <ENTRY entrytime="00:00:29.81" eventid="1133" heatid="40074" lane="8">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:29.81" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.26" eventid="1173" heatid="40139" lane="1">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:29.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.24" eventid="1237" heatid="40229" lane="7">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:08.83" />
                </ENTRY>
                <ENTRY entrytime="00:04:53.65" eventid="1257" heatid="40255" lane="2">
                  <MEETINFO name="Stadtwerke Erding Cup" city="Erding" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:04:50.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.42" eventid="1297" heatid="40335" lane="8" />
                <ENTRY entrytime="00:02:36.49" eventid="1317" heatid="40371" lane="4">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-11" qualificationtime="00:02:34.19" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.13" eventid="1357" heatid="40432" lane="7">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:17.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.21" eventid="1397" heatid="40491" lane="8">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:01:11.49" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Kaminski" birthdate="2012-01-01" gender="F" nation="GER" license="448677" athleteid="34726">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.36" eventid="1123" heatid="40037" lane="3">
                  <MEETINFO name="Bezirksmeisterschaften" city="Bobingen" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:32.36" />
                </ENTRY>
                <ENTRY entrytime="00:03:19.45" eventid="1143" heatid="40093" lane="8">
                  <MEETINFO name="38. Zirbelnuss-Schwimmen  des SV Augsburg 1911" city="Augsburg" course="SCM" approved="GER" date="2025-01-11" qualificationtime="00:03:19.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.01" eventid="1207" heatid="40165" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften" city="Bobingen" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:41.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.81" eventid="1227" heatid="40195" lane="4">
                  <MEETINFO name="Stadtberger Mehrkampftag" city="Stadtbergen" course="SCM" approved="GER" date="2025-04-27" qualificationtime="00:01:27.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.76" eventid="1267" heatid="40269" lane="6">
                  <MEETINFO name="Bezirksmeisterschaften" city="Bobingen" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:01:12.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.10" eventid="1327" heatid="40383" lane="2">
                  <MEETINFO name="Bezirksmeisterschaften" city="Bobingen" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:30.10" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.66" eventid="1347" heatid="40406" lane="5">
                  <MEETINFO name="Stadtberger Mehrkampftag" city="Stadtbergen" course="SCM" approved="GER" date="2025-04-27" qualificationtime="00:02:48.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.05" eventid="1367" heatid="40442" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Dornbusch" birthdate="2013-01-01" gender="M" nation="GER" license="448670" athleteid="34696">
              <ENTRIES>
                <ENTRY entrytime="00:20:51.14" eventid="1113" heatid="40023" lane="4">
                  <MEETINFO name="Bezirksmeistermeisterschaften Lange Strecke" city="Augsburg" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:19:39.39" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.82" eventid="1153" heatid="40106" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:56.43" />
                </ENTRY>
                <ENTRY entrytime="00:02:46.13" eventid="1173" heatid="40135" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:41.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.07" eventid="1217" heatid="40181" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:36.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.17" eventid="1237" heatid="40223" lane="7">
                  <MEETINFO name="Regionale Bestenkämpfe - Nord" city="Augsburg" course="SCM" approved="GER" date="2025-03-15" qualificationtime="00:01:15.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.83" eventid="1277" heatid="40297" lane="3">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:01:07.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.17" eventid="1337" heatid="40397" lane="7">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:19.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.25" eventid="1357" heatid="40428" lane="1">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:25.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.22" eventid="1377" heatid="40466" lane="6">
                  <MEETINFO name="2. SUN-SWIM Trophy" city="Neckarsulm" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:00:36.22" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:34.92" eventid="1185" heatid="40145" lane="6">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" date="2025-05-10" qualificationtime="00:01:55.14" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:35.66" eventid="1183" heatid="40143" lane="6">
                  <MEETINFO name="Bezirks-Jahrgangsmeisterschaften und Masters" city="Augsburg" date="2025-05-10" qualificationtime="00:02:13.66" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Christine" gender="M" lastname="Lienhart" />
            <COACH firstname="Christine" gender="M" lastname="Lienhart" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="0000" nation="CZE" clubid="35843" name="Plavecký klub Vodní stavby Praha">
          <CONTACT city="Prague" email="vosp@plavecky.club" internet="https://plavecky.club/" name="Michal Cervinka" state="CZE" />
          <ATHLETES>
            <ATHLETE firstname="Simon" lastname="Soban" birthdate="2011-05-26" gender="M" nation="CZE" athleteid="36371">
              <ENTRIES>
                <ENTRY entrytime="00:09:44.54" entrycourse="SCM" eventid="1093" heatid="40017" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:27.71" entrycourse="SCM" eventid="1133" heatid="40080" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:01:12.16" entrycourse="SCM" eventid="1237" heatid="40227" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:04:36.48" entrycourse="SCM" eventid="1257" heatid="40258" lane="2">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Florian" lastname="Fibir" birthdate="2011-02-16" gender="M" nation="CZE" athleteid="36332">
              <ENTRIES>
                <ENTRY entrytime="00:05:23.73" entrycourse="SCM" eventid="1073" heatid="40000" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:27.40" entrycourse="SCM" eventid="1133" heatid="40081" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:38.45" entrycourse="LCM" eventid="1217" heatid="40181" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:00.88" entrycourse="SCM" eventid="1277" heatid="40304" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:31.25" entrycourse="SCM" eventid="1297" heatid="40339" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:07.91" entrycourse="SCM" eventid="1397" heatid="40493" lane="8">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Barbora" lastname="Kacalova" birthdate="2010-08-12" gender="F" nation="CZE" athleteid="36357">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.77" entrycourse="SCM" eventid="1123" heatid="40042" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:03:00.50" entrycourse="SCM" eventid="1143" heatid="40097" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:00:39.22" entrycourse="SCM" eventid="1207" heatid="40168" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:01:09.10" entrycourse="SCM" eventid="1267" heatid="40275" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:00:35.22" entrycourse="SCM" eventid="1287" heatid="40317" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:25.15" entrycourse="SCM" eventid="1327" heatid="40387" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:00:40.79" entrycourse="LCM" eventid="1367" heatid="40442" lane="7">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sofie" lastname="Spurna" birthdate="2010-04-01" gender="F" nation="CZE" athleteid="36365">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.32" entrycourse="SCM" eventid="1123" heatid="40037" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:00:40.38" entrycourse="SCM" eventid="1207" heatid="40166" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:01:24.30" entrycourse="SCM" eventid="1227" heatid="40198" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:35.67" entrycourse="SCM" eventid="1287" heatid="40317" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:00:37.38" entrycourse="SCM" eventid="1367" heatid="40448" lane="3">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Fornusek" birthdate="2012-10-20" gender="M" nation="CZE" athleteid="36339">
              <ENTRIES>
                <ENTRY entrytime="00:19:38.00" entrycourse="SCM" eventid="1113" heatid="40024" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:38.33" entrycourse="SCM" eventid="1173" heatid="40137" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:01:15.01" entrycourse="SCM" eventid="1237" heatid="40225" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:06.81" entrycourse="SCM" eventid="1277" heatid="40298" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:44.09" entrycourse="SCM" eventid="1317" heatid="40370" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:02:24.24" entrycourse="SCM" eventid="1357" heatid="40429" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:00:35.51" entrycourse="SCM" eventid="1377" heatid="40467" lane="2">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maya" lastname="Haskova" birthdate="2013-04-17" gender="F" nation="CZE" athleteid="36347">
              <ENTRIES>
                <ENTRY entrytime="00:11:29.75" entrycourse="SCM" eventid="1083" heatid="40005" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:00:31.92" entrycourse="SCM" eventid="1123" heatid="40040" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:03:13.03" entrycourse="SCM" eventid="1143" heatid="40094" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:00:41.77" entrycourse="SCM" eventid="1207" heatid="40163" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:05:25.86" entrycourse="SCM" eventid="1247" heatid="40238" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:12.53" entrycourse="SCM" eventid="1267" heatid="40270" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:28.99" entrycourse="SCM" eventid="1327" heatid="40384" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:30.61" entrycourse="SCM" eventid="1347" heatid="40413" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:01:31.84" entrycourse="SCM" eventid="1387" heatid="40476" lane="4">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5555" nation="GER" region="16" clubid="36895" name="Erfurter SSC">
          <ATHLETES>
            <ATHLETE firstname="Sarafina" lastname="Schellhammer" birthdate="2012-01-01" gender="F" nation="GER" license="444321" athleteid="38474">
              <ENTRIES>
                <ENTRY entrytime="00:10:45.00" eventid="1083" heatid="40008" lane="4" />
                <ENTRY entrytime="00:00:30.95" eventid="1123" heatid="40046" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:31.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.67" eventid="1163" heatid="40124" lane="6">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:02:39.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.69" eventid="1207" heatid="40165" lane="3">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:40.69" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.75" eventid="1227" heatid="40209" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:13.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.40" eventid="1267" heatid="40277" lane="8">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:07.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.50" eventid="1287" heatid="40322" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:33.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.72" eventid="1367" heatid="40456" lane="6">
                  <MEETINFO name="Jugend trainert für Olympia" city="Berlin" course="SCM" approved="GER" date="2025-09-23" qualificationtime="00:00:33.60" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Florian" lastname="Eichelkraut" birthdate="2009-01-01" gender="M" nation="GER" license="382374" athleteid="38471">
              <ENTRIES>
                <ENTRY entrytime="00:02:23.76" eventid="1173" heatid="40140" lane="1">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:17.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.65" eventid="1197" heatid="40155" lane="3">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:17.40" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3266" nation="GER" region="16" clubid="34142" name="Meininger SV &quot;Wasserfreunde&quot; e.V.">
          <ATHLETES>
            <ATHLETE firstname="Moritz" lastname="Göpfert" birthdate="2013-01-01" gender="M" nation="GER" license="446198" athleteid="34143">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.87" eventid="1133" heatid="40062" lane="1">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:34.26" />
                </ENTRY>
                <ENTRY entrytime="00:03:15.90" eventid="1173" heatid="40129" lane="2">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:03:07.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.99" eventid="1237" heatid="40216" lane="5">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:01:29.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.54" eventid="1277" heatid="40290" lane="8">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:16.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.09" eventid="1357" heatid="40422" lane="3">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:54.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Luke" lastname="Reckwell" birthdate="2014-01-01" gender="M" nation="GER" license="446203" athleteid="34163">
              <ENTRIES>
                <ENTRY entrytime="00:03:29.01" eventid="1153" heatid="40103" lane="1">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:03:27.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.80" eventid="1237" heatid="40217" lane="2">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:26.45" />
                </ENTRY>
                <ENTRY entrytime="00:03:09.21" eventid="1317" heatid="40364" lane="2">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-26" qualificationtime="00:03:02.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.85" eventid="1357" heatid="40422" lane="4">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:48.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:42.21" eventid="1397" heatid="40486" lane="4">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:01:41.98" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anni" lastname="Reiß" birthdate="2015-01-01" gender="F" nation="GER" license="459776" athleteid="34169">
              <ENTRIES>
                <ENTRY entrytime="00:03:24.46" eventid="1163" heatid="40113" lane="8">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:03:19.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.27" eventid="1227" heatid="40193" lane="6">
                  <MEETINFO name="33. Internationale Geraer Stadtmeisterschaften" city="Gera" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:34.27" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.11" eventid="1267" heatid="40262" lane="3">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:01:20.37" />
                </ENTRY>
                <ENTRY entrytime="00:03:26.73" eventid="1307" heatid="40348" lane="5">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:03:21.98" />
                </ENTRY>
                <ENTRY entrytime="00:03:02.10" eventid="1347" heatid="40405" lane="2">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:50.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:48.53" eventid="1387" heatid="40475" lane="5">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:01:42.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Hoffmann" birthdate="2015-01-01" gender="M" nation="GER" license="465140" athleteid="34149">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.84" eventid="1133" heatid="40065" lane="8">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-26" qualificationtime="00:00:33.64" />
                </ENTRY>
                <ENTRY entrytime="00:03:23.22" eventid="1173" heatid="40128" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:03:08.90" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.99" eventid="1237" heatid="40216" lane="4">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:01:29.36" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.98" eventid="1277" heatid="40291" lane="1">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:16.84" />
                </ENTRY>
                <ENTRY entrytime="00:03:13.48" eventid="1317" heatid="40363" lane="3">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:03:01.49" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.04" eventid="1397" heatid="40487" lane="8">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:01:33.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fynn Leandro" lastname="Marr" birthdate="2014-01-01" gender="M" nation="GER" license="461903" athleteid="34156">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.87" eventid="1133" heatid="40061" lane="1">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:35.03" />
                </ENTRY>
                <ENTRY entrytime="00:03:21.05" eventid="1173" heatid="40128" lane="3">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:03:02.16" />
                </ENTRY>
                <ENTRY entrytime="00:05:48.14" eventid="1257" heatid="40248" lane="8">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:05:52.08" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.62" eventid="1277" heatid="40290" lane="5">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:01:17.72" />
                </ENTRY>
                <ENTRY entrytime="00:03:14.14" eventid="1317" heatid="40363" lane="6">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-26" qualificationtime="00:03:08.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.75" eventid="1397" heatid="40487" lane="4">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-25" qualificationtime="00:01:34.09" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Steiner" birthdate="2012-01-01" gender="M" nation="GER" license="446207" athleteid="34176">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.12" eventid="1133" heatid="40066" lane="5">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-26" qualificationtime="00:00:30.97" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.14" eventid="1173" heatid="40130" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:02:50.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.78" eventid="1217" heatid="40179" lane="7">
                  <MEETINFO name="Offene Thüringer Meisterschaften" city="Erfurt" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:00:40.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.14" eventid="1297" heatid="40334" lane="1">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-26" qualificationtime="00:00:35.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.32" eventid="1337" heatid="40396" lane="3">
                  <MEETINFO name="Thüringer Mehrkampfpokal und KIDS-CUP" city="Arnstadt" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:01:28.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.69" eventid="1397" heatid="40489" lane="2">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:17.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Jörg" gender="M" lastname="Kleinsteiber" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="4163" nation="GER" region="02" clubid="34817" name="1.FCN Schwimmen">
          <ATHLETES>
            <ATHLETE firstname="Fabian" lastname="Knorr" birthdate="2007-01-01" gender="M" nation="GER" license="377901" athleteid="35594">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.44" eventid="1133" heatid="40087" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:24.73" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.88" eventid="1153" heatid="40107" lane="4" />
                <ENTRY entrytime="00:00:31.40" eventid="1217" heatid="40189" lane="8">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:00:31.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.69" eventid="1277" heatid="40310" lane="8">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:54.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.94" eventid="1297" heatid="40345" lane="8">
                  <MEETINFO name="Offene Thüringer Meisterschaften" city="Erfurt" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:27.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.14" eventid="1337" heatid="40401" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:10.73" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.08" eventid="1357" heatid="40436" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Segerer" birthdate="2005-01-01" gender="F" nation="GER" license="368182" athleteid="35610">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.66" eventid="1123" heatid="40047" lane="3">
                  <MEETINFO name="Kreismeisterschaften Nord-Ost Mittelfranken" city="Lauf" course="SCM" approved="GER" date="2025-01-25" qualificationtime="00:00:30.02" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.19" eventid="1163" heatid="40120" lane="6">
                  <MEETINFO name="Kreismeisterschaften Nord-Ost Mittelfranken" city="Lauf" course="SCM" approved="GER" date="2025-01-25" qualificationtime="00:02:47.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.47" eventid="1207" heatid="40167" lane="3">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:39.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.07" eventid="1227" heatid="40204" lane="6">
                  <MEETINFO name="Int. Bayerische Kurzbahnmeisterschaften Masters" city="Fürstenfeldbruck" course="SCM" approved="GER" date="2025-03-22" qualificationtime="00:01:15.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.73" eventid="1267" heatid="40277" lane="4">
                  <MEETINFO name="Kreismeisterschaften Nord-Ost Mittelfranken" city="Lauf" course="SCM" approved="GER" date="2025-01-25" qualificationtime="00:01:07.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.44" eventid="1287" heatid="40319" lane="5">
                  <MEETINFO name="Bezirks- Jahrgangs- und Juniorenmeisterschaft KB" city="Nürnberg" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:34.44" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.97" eventid="1307" heatid="40357" lane="2">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:02:52.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.71" eventid="1367" heatid="40451" lane="5">
                  <MEETINFO name="Bezirks- Jahrgangs- und Juniorenmeisterschaft KB" city="Nürnberg" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:34.82" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Robin" lastname="Lienhart" birthdate="2006-01-01" gender="M" nation="GER" license="349208" athleteid="35602">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.53" eventid="1133" heatid="40088" lane="5">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:23.81" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.36" eventid="1153" heatid="40111" lane="2">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:02:16.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.71" eventid="1197" heatid="40156" lane="5">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-13" qualificationtime="00:02:02.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.26" eventid="1277" heatid="40311" lane="2">
                  <MEETINFO name="38. Zirbelnuss-Schwimmen  des SV Augsburg 1911" city="Augsburg" course="SCM" approved="GER" date="2025-01-12" qualificationtime="00:00:51.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.83" eventid="1297" heatid="40347" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:25.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.87" eventid="1337" heatid="40403" lane="7">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-13" qualificationtime="00:01:02.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.25" eventid="1397" heatid="40497" lane="1">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:55.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Jochen" gender="M" lastname="Stetina" />
            <COACH firstname="Julius" gender="M" lastname="Schönheid" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="3366" nation="GER" region="12" clubid="37970" name="SV Weixdorf e.V.">
          <ATHLETES>
            <ATHLETE firstname="Finja" lastname="Seidel" birthdate="2008-01-01" gender="F" nation="GER" license="349387" athleteid="37971">
              <ENTRIES>
                <ENTRY entrytime="00:17:36.86" eventid="1103" heatid="40021" lane="4">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:17:54.68" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.63" eventid="1143" heatid="40099" lane="8">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:02:48.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.44" eventid="1163" heatid="40127" lane="8">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:02:31.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.47" eventid="1227" heatid="40213" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:08.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.41" eventid="1307" heatid="40360" lane="6">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:02:31.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.32" eventid="1327" heatid="40390" lane="8">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:20.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Albrecht" birthdate="2010-01-01" gender="F" nation="GER" license="404147" athleteid="37978">
              <ENTRIES>
                <ENTRY entrytime="00:09:20.36" eventid="1083" heatid="40011" lane="5">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:09:20.36" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.02" eventid="1187" heatid="40150" lane="5">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:02:22.02" />
                </ENTRY>
                <ENTRY entrytime="00:04:25.72" eventid="1247" heatid="40245" lane="5">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:04:25.72" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.08" eventid="1347" heatid="40420" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:09.50" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Dorothea" lastname="Koenig" birthdate="2013-01-01" gender="F" nation="GER" license="424080" athleteid="37983">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.42" eventid="1123" heatid="40053" lane="7">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:29.42" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.43" eventid="1163" heatid="40122" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:40.17" />
                </ENTRY>
                <ENTRY entrytime="00:05:29.27" eventid="1247" heatid="40237" lane="4" />
                <ENTRY entrytime="00:02:52.28" eventid="1307" heatid="40355" lane="2" />
                <ENTRY entrytime="00:02:25.22" eventid="1347" heatid="40416" lane="3">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:02:25.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.01" eventid="1367" heatid="40455" lane="6">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:32.78" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Koenig" birthdate="2007-01-01" gender="M" nation="GER" license="333012" athleteid="37990">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.97" eventid="1133" heatid="40086" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:25.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.90" eventid="1277" heatid="40309" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:56.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.65" eventid="1297" heatid="40345" lane="1">
                  <MEETINFO name="Int. BAUAkademie ATUS Graz Trophy" city="Graz" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:00:27.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6524" nation="GER" region="02" clubid="34278" name="SC Regensburg">
          <ATHLETES>
            <ATHLETE firstname="Maya Zoe" lastname="Orth" birthdate="2011-01-01" gender="F" nation="GER" license="424437" athleteid="36141">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.82" eventid="1123" heatid="40051" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:29.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:46.82" eventid="1163" heatid="40121" lane="2">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:43.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.08" eventid="1227" heatid="40207" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:15.58" />
                </ENTRY>
                <ENTRY entrytime="00:05:09.20" eventid="1247" heatid="40242" lane="6">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:05:11.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.67" eventid="1267" heatid="40280" lane="2">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:05.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.98" eventid="1287" heatid="40321" lane="1">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:32.54" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.77" eventid="1307" heatid="40354" lane="3">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:53.77" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alexander" lastname="Hutchinson Riquelme" birthdate="2013-01-01" gender="M" nation="GER" license="443849" athleteid="36030">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.56" eventid="1133" heatid="40063" lane="4">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:34.25" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.26" eventid="1173" heatid="40131" lane="1">
                  <MEETINFO name="XVIII Meeting di Nuoto" city="Lignano Sabbiadoro" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:03:01.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.76" eventid="1237" heatid="40218" lane="3">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:23.46" />
                </ENTRY>
                <ENTRY entrytime="00:05:31.79" eventid="1257" heatid="40249" lane="7">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:05:26.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.98" eventid="1297" heatid="40336" lane="2">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:33.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.65" eventid="1317" heatid="40368" lane="6">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:48.60" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.84" eventid="1357" heatid="40425" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:32.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.71" eventid="1377" heatid="40462" lane="8">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:40.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Szemen" lastname="Matyuhin" birthdate="2011-01-01" gender="M" nation="GER" license="423598" athleteid="36068">
              <ENTRIES>
                <ENTRY entrytime="00:19:00.99" eventid="1113" heatid="40025" lane="1">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-10" qualificationtime="00:19:20.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.50" eventid="1133" heatid="40077" lane="4">
                  <MEETINFO name="Kreisjahrgangsmeisterschaften Ost" city="Viechtach" course="SCM" approved="GER" date="2025-02-22" qualificationtime="00:00:27.41" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.99" eventid="1153" heatid="40109" lane="4">
                  <MEETINFO name="Niederbayerische Langbahnmeisterschaften" city="Mainburg" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:40.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.59" eventid="1217" heatid="40188" lane="1">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:32.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.99" eventid="1277" heatid="40304" lane="7">
                  <MEETINFO name="Kreisjahrgangsmeisterschaften Ost" city="Viechtach" course="SCM" approved="GER" date="2025-02-22" qualificationtime="00:00:59.79" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.99" eventid="1337" heatid="40402" lane="8">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:10.60" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Schaffarzik" birthdate="2011-01-01" gender="F" nation="GER" license="476624" athleteid="36204">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.99" eventid="1123" heatid="40039" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:30.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.50" eventid="1207" heatid="40162" lane="6">
                  <MEETINFO name="6. CabrioSol Cup Pegnitz" city="Pegnitz" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:42.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.00" eventid="1287" heatid="40320" lane="5">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:33.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.99" eventid="1307" heatid="40353" lane="3" />
                <ENTRY entrytime="00:01:28.99" eventid="1327" heatid="40384" lane="6" />
                <ENTRY entrytime="00:00:37.50" eventid="1367" heatid="40448" lane="2">
                  <MEETINFO name="6. CabrioSol Cup Pegnitz" city="Pegnitz" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:36.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.99" eventid="1387" heatid="40479" lane="2">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:24.34" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jacob" lastname="Mulzer" birthdate="2014-01-01" gender="M" nation="GER" license="449265" athleteid="36084">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.19" eventid="1133" heatid="40060" lane="5">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:00:37.19" />
                </ENTRY>
                <ENTRY entrytime="00:03:17.83" eventid="1173" heatid="40129" lane="1">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:03:17.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.00" eventid="1237" heatid="40215" lane="2">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:31.15" />
                </ENTRY>
                <ENTRY entrytime="00:05:55.00" eventid="1257" heatid="40247" lane="6">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:05:58.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.30" eventid="1277" heatid="40288" lane="3">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:17.63" />
                </ENTRY>
                <ENTRY entrytime="00:03:16.12" eventid="1317" heatid="40363" lane="1">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:03:06.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.33" eventid="1357" heatid="40423" lane="1">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:47.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.84" eventid="1377" heatid="40461" lane="2">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:43.84" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Linda" lastname="Mahl" birthdate="2013-01-01" gender="F" nation="GER" license="443844" athleteid="36049">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.16" eventid="1123" heatid="40032" lane="1">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:33.25" />
                </ENTRY>
                <ENTRY entrytime="00:03:09.34" eventid="1143" heatid="40094" lane="5">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:03:09.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.86" eventid="1207" heatid="40165" lane="2">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:40.86" />
                </ENTRY>
                <ENTRY entrytime="00:05:36.45" eventid="1247" heatid="40237" lane="7">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:05:36.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.75" eventid="1287" heatid="40315" lane="8">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-17" qualificationtime="00:00:36.75" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.09" eventid="1307" heatid="40353" lane="6">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:49.49" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.34" eventid="1327" heatid="40385" lane="3">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:27.28" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.26" eventid="1347" heatid="40410" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:36.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.00" eventid="1367" heatid="40444" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Amira" lastname="Varna" birthdate="2006-01-01" gender="F" nation="GER" license="358238" athleteid="36280">
              <ENTRIES>
                <ENTRY entrytime="00:02:35.99" eventid="1163" heatid="40125" lane="3" />
                <ENTRY entrytime="00:01:10.93" eventid="1227" heatid="40211" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:08.93" />
                </ENTRY>
                <ENTRY entrytime="00:04:42.98" eventid="1247" heatid="40245" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:04:38.98" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.05" eventid="1267" heatid="40283" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:01.04" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.21" eventid="1347" heatid="40419" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:13.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Klara" lastname="Nagler" birthdate="2012-01-01" gender="F" nation="GER" license="442816" athleteid="36112">
              <ENTRIES>
                <ENTRY entrytime="00:06:02.77" eventid="1063" heatid="39995" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:05:51.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.40" eventid="1123" heatid="40037" lane="2">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:32.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.03" eventid="1163" heatid="40119" lane="6">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:50.03" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.18" eventid="1187" heatid="40150" lane="8">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:02:39.18" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.37" eventid="1227" heatid="40202" lane="1">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:18.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.64" eventid="1267" heatid="40269" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:10.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.95" eventid="1287" heatid="40323" lane="4">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:32.95" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.31" eventid="1307" heatid="40356" lane="4">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:02:47.31" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.11" eventid="1347" heatid="40411" lane="1">
                  <MEETINFO name="Kleines Märzmeeting" city="Nürnberg" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:37.11" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.02" eventid="1387" heatid="40483" lane="6">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:01:12.02" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Andrew" lastname="Cicero" birthdate="2010-01-01" gender="M" nation="GER" license="412140" athleteid="35990">
              <ENTRIES>
                <ENTRY entrytime="00:09:39.19" eventid="1093" heatid="40017" lane="5">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:09:22.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.37" eventid="1133" heatid="40078" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:27.19" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.56" eventid="1173" heatid="40140" lane="7">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:02:23.56" />
                </ENTRY>
                <ENTRY entrytime="00:04:23.70" eventid="1257" heatid="40259" lane="2">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:04:16.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.41" eventid="1277" heatid="40307" lane="1">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:57.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.04" eventid="1297" heatid="40340" lane="2">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-12" qualificationtime="00:00:31.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.59" eventid="1357" heatid="40437" lane="7">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:02.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.10" eventid="1377" heatid="40471" lane="7">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:29.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Rebeka" lastname="Voznak" birthdate="2015-01-01" gender="F" nation="GER" license="464352" athleteid="36286">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.54" eventid="1123" heatid="40043" lane="6">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:00:31.54" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.86" eventid="1163" heatid="40115" lane="8">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:03:05.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.00" eventid="1227" heatid="40197" lane="5">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:26.08" />
                </ENTRY>
                <ENTRY entrytime="00:05:44.92" eventid="1247" heatid="40236" lane="2">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-18" qualificationtime="00:05:44.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.45" eventid="1287" heatid="40319" lane="3">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:34.45" />
                </ENTRY>
                <ENTRY entrytime="00:03:02.41" eventid="1307" heatid="40351" lane="5">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:03:02.41" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.04" eventid="1347" heatid="40408" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:41.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.78" eventid="1367" heatid="40445" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:38.78" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jovana" lastname="Todorovska" birthdate="2014-01-01" gender="F" nation="MKD" license="478503" athleteid="36257">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.93" eventid="1123" heatid="40046" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:29.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.10" eventid="1163" heatid="40123" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:36.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.16" eventid="1227" heatid="40209" lane="6">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:01:10.06" />
                </ENTRY>
                <ENTRY entrytime="00:05:09.79" eventid="1247" heatid="40242" lane="2">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-18" qualificationtime="00:05:09.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.45" eventid="1287" heatid="40325" lane="2">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:31.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.24" eventid="1307" heatid="40357" lane="6">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:36.26" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.34" eventid="1347" heatid="40416" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:24.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.58" eventid="1367" heatid="40454" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:32.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Johanna Malene" lastname="Hecht" birthdate="2014-01-01" gender="F" nation="GER" license="455010" athleteid="36015">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.45" eventid="1123" heatid="40034" lane="7">
                  <MEETINFO name="Niederbayerische Langbahnmeisterschaften" city="Mainburg" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:33.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.81" eventid="1163" heatid="40118" lane="4">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:02:51.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.61" eventid="1207" heatid="40158" lane="2">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:46.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.19" eventid="1227" heatid="40205" lane="7">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:17.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Louisa" lastname="Muñoz" birthdate="2014-01-01" gender="F" nation="GER" license="457808" athleteid="36093">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.54" eventid="1123" heatid="40027" lane="4">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:36.54" />
                </ENTRY>
                <ENTRY entrytime="00:03:45.00" eventid="1143" heatid="40090" lane="1">
                  <MEETINFO name="International Swim Meeting" city="Erlangen" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:03:56.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.61" eventid="1227" heatid="40196" lane="3">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:26.61" />
                </ENTRY>
                <ENTRY entrytime="00:05:55.00" eventid="1247" heatid="40235" lane="2">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:06:10.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.81" eventid="1287" heatid="40313" lane="3">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:38.81" />
                </ENTRY>
                <ENTRY entrytime="00:03:12.82" eventid="1307" heatid="40349" lane="2">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:03:05.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:49.47" eventid="1327" heatid="40378" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:46.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:57.61" eventid="1347" heatid="40406" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:55.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.29" eventid="1367" heatid="40441" lane="8">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:42.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Damjan" lastname="Todorovski" birthdate="2009-01-01" gender="M" nation="MKD" license="478502" athleteid="36266">
              <ENTRIES>
                <ENTRY entrytime="00:02:34.76" eventid="1153" heatid="40110" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:02:34.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.73" eventid="1217" heatid="40189" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:29.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.80" eventid="1237" heatid="40227" lane="1">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:12.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.65" eventid="1297" heatid="40342" lane="2">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:29.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.34" eventid="1337" heatid="40402" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:06.35" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.21" eventid="1357" heatid="40434" lane="1">
                  <MEETINFO name="XVIII Meeting di Nuoto" city="Lignano Sabbiadoro" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:02:13.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Rummel" birthdate="2014-01-01" gender="F" nation="GER" license="458196" athleteid="36193">
              <ENTRIES>
                <ENTRY entrytime="00:11:30.00" eventid="1083" heatid="40005" lane="1" />
                <ENTRY entrytime="00:03:24.20" eventid="1143" heatid="40092" lane="7">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:03:24.20" />
                </ENTRY>
                <ENTRY entrytime="00:03:10.38" eventid="1163" heatid="40114" lane="8">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:03:10.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.34" eventid="1207" heatid="40158" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:00:45.78" />
                </ENTRY>
                <ENTRY entrytime="00:05:39.05" eventid="1247" heatid="40236" lane="5">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-18" qualificationtime="00:05:39.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.13" eventid="1267" heatid="40266" lane="2">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:16.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.27" eventid="1307" heatid="40352" lane="2">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:02:58.27" />
                </ENTRY>
                <ENTRY entrytime="00:01:38.59" eventid="1327" heatid="40380" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:35.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.16" eventid="1347" heatid="40408" lane="7">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:44.16" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.98" eventid="1367" heatid="40440" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:43.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Greta" lastname="Oberneder" birthdate="2012-01-01" gender="F" nation="GER" license="458074" athleteid="36133">
              <ENTRIES>
                <ENTRY entrytime="00:05:45.99" eventid="1063" heatid="39996" lane="2" />
                <ENTRY entrytime="00:02:50.99" eventid="1163" heatid="40119" lane="7">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:02:54.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.74" eventid="1227" heatid="40201" lane="3">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:18.11" />
                </ENTRY>
                <ENTRY entrytime="00:05:20.99" eventid="1247" heatid="40239" lane="8" />
                <ENTRY entrytime="00:00:32.99" eventid="1287" heatid="40323" lane="3">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:00:32.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.12" eventid="1307" heatid="40354" lane="2">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:47.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.02" eventid="1387" heatid="40482" lane="4">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:14.02" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Mahl" birthdate="2010-01-01" gender="F" nation="GER" license="414341" athleteid="36059">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.63" eventid="1123" heatid="40052" lane="8">
                  <MEETINFO name="Kleines Märzmeeting" city="Nürnberg" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:29.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.21" eventid="1163" heatid="40121" lane="5">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:38.16" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.82" eventid="1227" heatid="40206" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:13.41" />
                </ENTRY>
                <ENTRY entrytime="00:04:55.99" eventid="1247" heatid="40243" lane="6">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:04:59.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.92" eventid="1267" heatid="40281" lane="6">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:04.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.11" eventid="1287" heatid="40320" lane="3">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:00:34.34" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.39" eventid="1347" heatid="40417" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:17.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.60" eventid="1367" heatid="40454" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:33.22" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Stangelmayer" birthdate="2010-01-01" gender="F" nation="GER" license="414346" athleteid="36240">
              <ENTRIES>
                <ENTRY entrytime="00:02:56.92" eventid="1143" heatid="40098" lane="7">
                  <MEETINFO name="2. Nürnberger Schwimmfest" city="Nürnberg" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:02:57.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.49" eventid="1207" heatid="40167" lane="2">
                  <MEETINFO name="Kleines Märzmeeting" city="Nürnberg" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:39.49" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.72" eventid="1227" heatid="40199" lane="7" />
                <ENTRY entrytime="00:01:07.42" eventid="1267" heatid="40278" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:07.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.48" eventid="1287" heatid="40322" lane="1">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-17" qualificationtime="00:00:33.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.79" eventid="1327" heatid="40388" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:22.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.64" eventid="1367" heatid="40448" lane="8">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:36.44" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Nowey" birthdate="2013-01-01" gender="M" nation="GER" license="443841" athleteid="36123">
              <ENTRIES>
                <ENTRY entrytime="00:02:51.53" eventid="1153" heatid="40108" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:45.81" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.31" eventid="1173" heatid="40130" lane="4">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:03:03.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.94" eventid="1217" heatid="40182" lane="1">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:37.15" />
                </ENTRY>
                <ENTRY entrytime="00:05:36.26" eventid="1257" heatid="40249" lane="8">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:05:19.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.70" eventid="1297" heatid="40333" lane="5">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:00:35.38" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.86" eventid="1317" heatid="40368" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:40.38" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.54" eventid="1337" heatid="40398" lane="1">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:18.28" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.25" eventid="1357" heatid="40426" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:28.90" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.85" eventid="1377" heatid="40463" lane="6">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:39.85" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maxim" lastname="Belyaev" birthdate="2012-01-01" gender="M" nation="GER" license="442808" athleteid="35979">
              <ENTRIES>
                <ENTRY entrytime="00:05:45.52" eventid="1073" heatid="40000" lane="8">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-12" qualificationtime="00:06:07.52" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.98" eventid="1133" heatid="40073" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:28.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.02" eventid="1173" heatid="40136" lane="7">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:02:42.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.59" eventid="1237" heatid="40225" lane="3">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:10.74" />
                </ENTRY>
                <ENTRY entrytime="00:05:02.42" eventid="1257" heatid="40254" lane="6">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:05:02.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.09" eventid="1277" heatid="40300" lane="4">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:01.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.56" eventid="1297" heatid="40334" lane="6">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:00:34.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.89" eventid="1317" heatid="40370" lane="2">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:43.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.00" eventid="1357" heatid="40430" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:19.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.46" eventid="1377" heatid="40467" lane="3">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:34.42" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Helene" lastname="Herdeg" birthdate="2012-01-01" gender="F" nation="GER" license="443834" athleteid="36020">
              <ENTRIES>
                <ENTRY entrytime="00:10:53.99" eventid="1083" heatid="40008" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:10:40.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.77" eventid="1123" heatid="40042" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:31.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.80" eventid="1227" heatid="40199" lane="1">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:23.80" />
                </ENTRY>
                <ENTRY entrytime="00:05:10.36" eventid="1247" heatid="40242" lane="1">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:05:10.36" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.26" eventid="1267" heatid="40274" lane="4">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-17" qualificationtime="00:01:09.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.02" eventid="1287" heatid="40316" lane="2">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:35.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.24" eventid="1307" heatid="40353" lane="5">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:50.25" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.96" eventid="1347" heatid="40415" lane="8">
                  <MEETINFO name="17. Intern Franz v. Kirchbauer Gedächtnisschwimmen" city="Burghausen" course="LCM" approved="GER" date="2025-05-17" qualificationtime="00:02:27.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.99" eventid="1387" heatid="40477" lane="4">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:21.54" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Kilian" lastname="Sußbauer" birthdate="2013-01-01" gender="M" nation="GER" license="445749" athleteid="36248">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.33" eventid="1133" heatid="40061" lane="5">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:36.29" />
                </ENTRY>
                <ENTRY entrytime="00:03:08.62" eventid="1173" heatid="40130" lane="7">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-12" qualificationtime="00:03:08.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.69" eventid="1237" heatid="40217" lane="5">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:24.08" />
                </ENTRY>
                <ENTRY entrytime="00:05:40.00" eventid="1257" heatid="40248" lane="6">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:06:09.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.57" eventid="1277" heatid="40289" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:17.80" />
                </ENTRY>
                <ENTRY entrytime="00:03:10.10" eventid="1317" heatid="40364" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:58.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.36" eventid="1357" heatid="40423" lane="8">
                  <MEETINFO name="XVIII Meeting di Nuoto" city="Lignano Sabbiadoro" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:02:53.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.52" eventid="1377" heatid="40462" lane="7">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:41.52" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emma" lastname="Irrgang" birthdate="2012-01-01" gender="F" nation="GER" license="443835" athleteid="36039">
              <ENTRIES>
                <ENTRY entrytime="00:10:04.10" eventid="1083" heatid="40010" lane="3">
                  <MEETINFO name="Bay. Meisterschaften Lange Strecken" city="Würzburg" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:10:04.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.42" eventid="1123" heatid="40053" lane="1">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:00:29.42" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.34" eventid="1163" heatid="40126" lane="6">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:31.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.78" eventid="1227" heatid="40211" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:10.59" />
                </ENTRY>
                <ENTRY entrytime="00:04:51.97" eventid="1247" heatid="40244" lane="1">
                  <MEETINFO name="Bay. Meisterschaften Lange Strecken" city="Würzburg" course="LCM" approved="GER" date="2025-01-18" qualificationtime="00:04:51.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.92" eventid="1267" heatid="40283" lane="5">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:01:02.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.16" eventid="1307" heatid="40359" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:02:32.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.07" eventid="1347" heatid="40419" lane="8">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:16.37" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.95" eventid="1387" heatid="40484" lane="7">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:01:10.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Julia Pia" lastname="Schüller" birthdate="2011-01-01" gender="F" nation="GER" license="443830" athleteid="36221">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.68" eventid="1123" heatid="40047" lane="2">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:00:30.68" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.95" eventid="1163" heatid="40117" lane="6" />
                <ENTRY entrytime="00:01:21.32" eventid="1227" heatid="40202" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:19.53" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.91" eventid="1247" heatid="40240" lane="2" />
                <ENTRY entrytime="00:01:09.41" eventid="1267" heatid="40274" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:09.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.91" eventid="1287" heatid="40321" lane="2">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-12" qualificationtime="00:00:33.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.67" eventid="1347" heatid="40410" lane="3" />
                <ENTRY entrytime="00:00:37.10" eventid="1367" heatid="40448" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:36.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Raúl" lastname="Muñoz" birthdate="2011-01-01" gender="M" nation="GER" license="424436" athleteid="36103">
              <ENTRIES>
                <ENTRY entrytime="00:10:10.00" eventid="1093" heatid="40016" lane="5">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:10:16.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.14" eventid="1133" heatid="40075" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:28.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.13" eventid="1173" heatid="40134" lane="8">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:02:51.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.92" eventid="1237" heatid="40223" lane="3">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:13.49" />
                </ENTRY>
                <ENTRY entrytime="00:04:42.95" eventid="1257" heatid="40257" lane="8">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-18" qualificationtime="00:04:42.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.23" eventid="1277" heatid="40303" lane="7">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:01:02.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.86" eventid="1357" heatid="40433" lane="7">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:02:14.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.23" eventid="1377" heatid="40466" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:35.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Osteroth" birthdate="2009-01-01" gender="F" nation="GER" license="400513" athleteid="36159">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.52" eventid="1123" heatid="40043" lane="3">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-12" qualificationtime="00:00:31.52" />
                </ENTRY>
                <ENTRY entrytime="00:03:06.54" eventid="1143" heatid="40095" lane="3" />
                <ENTRY entrytime="00:02:58.16" eventid="1187" heatid="40148" lane="2" />
                <ENTRY entrytime="00:00:38.43" eventid="1207" heatid="40169" lane="3">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-11" qualificationtime="00:00:38.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.66" eventid="1267" heatid="40272" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:07.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.73" eventid="1327" heatid="40386" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:26.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Gross" birthdate="2010-01-01" gender="M" nation="GER" license="415119" athleteid="36006">
              <ENTRIES>
                <ENTRY entrytime="00:05:20.98" eventid="1073" heatid="40000" lane="5">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:05:32.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.40" eventid="1133" heatid="40081" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:27.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.99" eventid="1197" heatid="40152" lane="6" />
                <ENTRY entrytime="00:01:12.16" eventid="1237" heatid="40227" lane="3">
                  <MEETINFO name="6. CabrioSol Cup Pegnitz" city="Pegnitz" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:11.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.60" eventid="1277" heatid="40306" lane="6">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:58.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.03" eventid="1317" heatid="40372" lane="7">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:02:35.03" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.37" eventid="1357" heatid="40434" lane="8">
                  <MEETINFO name="DMS-Austragung 24/25 Bezirksliga - Oberpfalz" city="Weiden" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:02:10.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.00" eventid="1397" heatid="40491" lane="1">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:08.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marc" lastname="Rohrmüller" birthdate="2011-01-01" gender="M" nation="GER" license="424439" athleteid="36174">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.59" eventid="1133" heatid="40080" lane="4">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:26.44" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.37" eventid="1197" heatid="40152" lane="4">
                  <MEETINFO name="DMS-Austragung 24/25 Bezirksliga - Oberpfalz" city="Weiden" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:02:52.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.97" eventid="1277" heatid="40307" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:57.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.94" eventid="1297" heatid="40343" lane="3">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:28.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.26" eventid="1357" heatid="40435" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:10.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.15" eventid="1397" heatid="40492" lane="8">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:06.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Ostermeier" birthdate="2012-01-01" gender="F" nation="GER" license="442817" athleteid="36149">
              <ENTRIES>
                <ENTRY entrytime="00:11:02.93" eventid="1083" heatid="40006" lane="4">
                  <MEETINFO name="Bay. Meisterschaften Lange Strecken" city="Würzburg" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:11:02.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.91" eventid="1123" heatid="40050" lane="6">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:00:29.91" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.66" eventid="1143" heatid="40096" lane="3">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:03:03.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.97" eventid="1207" heatid="40170" lane="5">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:00:37.97" />
                </ENTRY>
                <ENTRY entrytime="00:05:14.87" eventid="1247" heatid="40241" lane="1">
                  <MEETINFO name="XVIII Meeting di Nuoto" city="Lignano Sabbiadoro" course="LCM" approved="GER" date="2025-04-25" qualificationtime="00:05:14.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.09" eventid="1267" heatid="40281" lane="8">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:01:05.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.09" eventid="1307" heatid="40357" lane="4">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:02:43.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.42" eventid="1327" heatid="40386" lane="4">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:23.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.40" eventid="1347" heatid="40417" lane="5">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:22.40" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maximilian" lastname="Meier" birthdate="2013-01-01" gender="M" nation="GER" license="462715" athleteid="36075">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.61" eventid="1133" heatid="40065" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:32.72" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.19" eventid="1173" heatid="40132" lane="6">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:58.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.31" eventid="1237" heatid="40219" lane="2">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:24.30" />
                </ENTRY>
                <ENTRY entrytime="00:05:40.00" eventid="1257" heatid="40248" lane="3">
                  <MEETINFO name="Nürnberger Lange Strecken" city="Nürnberg" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:05:37.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.11" eventid="1277" heatid="40293" lane="4">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:13.01" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.87" eventid="1317" heatid="40366" lane="2">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:02:55.87" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.83" eventid="1357" heatid="40425" lane="6">
                  <MEETINFO name="XVIII Meeting di Nuoto" city="Lignano Sabbiadoro" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:02:36.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.05" eventid="1377" heatid="40463" lane="1">
                  <MEETINFO name="International Swim Meeting" city="Erlangen" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:40.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mia Luisa" lastname="Schönberger" birthdate="2011-01-01" gender="F" nation="GER" license="443832" athleteid="36212">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.80" eventid="1123" heatid="40042" lane="8">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:31.34" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.49" eventid="1163" heatid="40120" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:41.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.30" eventid="1227" heatid="40208" lane="7">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:11.40" />
                </ENTRY>
                <ENTRY entrytime="00:05:13.47" eventid="1247" heatid="40241" lane="6">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:05:13.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.28" eventid="1267" heatid="40274" lane="5">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:07.90" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.84" eventid="1327" heatid="40385" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:25.85" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.23" eventid="1347" heatid="40411" lane="2">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:36.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.37" eventid="1367" heatid="40455" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:33.45" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Dimitar" lastname="Todorovski" birthdate="2009-01-01" gender="M" nation="MKD" license="478501" athleteid="36273">
              <ENTRIES>
                <ENTRY entrytime="00:02:28.37" eventid="1153" heatid="40111" lane="7">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:24.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.49" eventid="1217" heatid="40189" lane="5">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:30.21" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.35" eventid="1237" heatid="40226" lane="7">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:14.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.69" eventid="1277" heatid="40308" lane="2">
                  <MEETINFO name="International Swim Meeting" city="Erlangen" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:59.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.04" eventid="1337" heatid="40402" lane="5">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:06.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.73" eventid="1357" heatid="40436" lane="1">
                  <MEETINFO name="XVIII Meeting di Nuoto" city="Lignano Sabbiadoro" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:02:08.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lina" lastname="Sinkel" birthdate="2011-01-01" gender="F" nation="GER" license="424441" athleteid="36230">
              <ENTRIES>
                <ENTRY entrytime="00:10:58.75" eventid="1083" heatid="40007" lane="4">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-10" qualificationtime="00:10:58.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.06" eventid="1123" heatid="40045" lane="3">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:31.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.65" eventid="1163" heatid="40120" lane="1">
                  <MEETINFO name="Swim Cup" city="Regensburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:49.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.37" eventid="1227" heatid="40203" lane="8">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:18.97" />
                </ENTRY>
                <ENTRY entrytime="00:05:10.40" eventid="1247" heatid="40242" lane="8">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-11" qualificationtime="00:05:16.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.20" eventid="1267" heatid="40277" lane="7">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:07.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.73" eventid="1287" heatid="40321" lane="6">
                  <MEETINFO name="29. Erlanger Röthelheimcup" city="Erlangen" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:00:33.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.96" eventid="1347" heatid="40414" lane="2">
                  <MEETINFO name="Kleines Märzmeeting" city="Nürnberg" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:28.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.05" eventid="1367" heatid="40449" lane="8">
                  <MEETINFO name="6. CabrioSol Cup Pegnitz" city="Pegnitz" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:36.83" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lia" lastname="Padberg" birthdate="2008-01-01" gender="F" nation="GER" license="390058" athleteid="36166">
              <ENTRIES>
                <ENTRY entrytime="00:10:00.53" eventid="1083" heatid="40010" lane="4">
                  <MEETINFO name="25. Internationaler Ratisbona-Cup" city="Regensburg" course="LCM" approved="GER" date="2025-01-10" qualificationtime="00:10:00.53" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.92" eventid="1163" heatid="40125" lane="4">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:32.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.80" eventid="1227" heatid="40210" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:11.59" />
                </ENTRY>
                <ENTRY entrytime="00:04:48.88" eventid="1247" heatid="40244" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:04:43.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.95" eventid="1267" heatid="40282" lane="5">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:03.75" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.25" eventid="1347" heatid="40419" lane="7">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:15.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.59" eventid="1367" heatid="40454" lane="2">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:33.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Franz" lastname="Rummel" birthdate="2011-01-01" gender="M" nation="GER" license="431792" athleteid="36181">
              <ENTRIES>
                <ENTRY entrytime="00:10:03.12" eventid="1093" heatid="40017" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:10:03.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.91" eventid="1133" heatid="40076" lane="3">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:28.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:46.82" eventid="1173" heatid="40135" lane="6">
                  <MEETINFO name="Sommermeisterschaften des Bezirks Oberpfalz" city="Weiden i. d. Opf." course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:02:46.82" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.97" eventid="1217" heatid="40182" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:37.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.92" eventid="1237" heatid="40225" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:14.72" />
                </ENTRY>
                <ENTRY entrytime="00:04:49.77" eventid="1257" heatid="40256" lane="8">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:04:49.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.32" eventid="1277" heatid="40301" lane="5">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:02.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.25" eventid="1317" heatid="40371" lane="2">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:37.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.43" eventid="1337" heatid="40397" lane="1">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:22.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.09" eventid="1357" heatid="40432" lane="6">
                  <MEETINFO name="Bezirkskurzbahnmeisterschaft Oberpfalz" city="Schwandorf" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:14.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.10" eventid="1377" heatid="40465" lane="2">
                  <MEETINFO name="Bayreuther Herbstme" city="Bayreuth" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:34.03" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Cicero" birthdate="2008-01-01" gender="M" nation="USA" license="412141" athleteid="35999">
              <ENTRIES>
                <ENTRY entrytime="00:08:45.50" eventid="1093" heatid="40019" lane="7" />
                <ENTRY entrytime="00:00:24.76" eventid="1133" heatid="40088" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:24.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.71" eventid="1237" heatid="40232" lane="4">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:53.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.58" eventid="1277" heatid="40311" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:53.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.23" eventid="1297" heatid="40347" lane="7">
                  <MEETINFO name="International Swim Meeting" city="Erlangen" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:26.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.17" eventid="1377" heatid="40474" lane="4">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:00:24.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:01:49.80" eventid="1185" heatid="40146" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="35999" number="1" />
                    <RELAYPOSITION athleteid="36266" number="2" />
                    <RELAYPOSITION athleteid="36174" number="3" />
                    <RELAYPOSITION athleteid="36273" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="24. Int. Dachauer Masters-Cup" city="Dachau" date="2025-02-22" qualificationtime="00:02:09.20" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.56" eventid="1185" heatid="40146" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="35990" number="1" />
                    <RELAYPOSITION athleteid="36068" number="2" />
                    <RELAYPOSITION athleteid="36006" number="3" />
                    <RELAYPOSITION athleteid="36181" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="24. Int. Dachauer Masters-Cup" city="Dachau" date="2025-02-22" qualificationtime="00:02:09.20" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <ENTRIES>
                <ENTRY entrytime="00:02:27.47" eventid="1185" heatid="40145" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="36075" number="1" />
                    <RELAYPOSITION athleteid="36123" number="2" />
                    <RELAYPOSITION athleteid="36030" number="3" />
                    <RELAYPOSITION athleteid="36248" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="24. Int. Dachauer Masters-Cup" city="Dachau" date="2025-02-22" qualificationtime="00:02:09.20" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:15.71" eventid="1183" heatid="40144" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="36039" number="1" />
                    <RELAYPOSITION athleteid="36240" number="2" />
                    <RELAYPOSITION athleteid="36280" number="3" />
                    <RELAYPOSITION athleteid="36059" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="15. Deutsche Kurzbahnmeisterschaft der Masters" city="Essen" date="2025-11-30" qualificationtime="00:02:10.88" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <ENTRIES>
                <ENTRY entrytime="00:02:14.66" eventid="1183" heatid="40144" lane="7">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="36166" number="1" />
                    <RELAYPOSITION athleteid="36159" number="2" />
                    <RELAYPOSITION athleteid="36112" number="3" />
                    <RELAYPOSITION athleteid="36149" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="15. Deutsche Kurzbahnmeisterschaft der Masters" city="Essen" date="2025-11-30" qualificationtime="00:02:10.88" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <ENTRIES>
                <ENTRY entrytime="00:02:21.57" eventid="1183" heatid="40143" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="36230" number="1" />
                    <RELAYPOSITION athleteid="36204" number="2" />
                    <RELAYPOSITION athleteid="36133" number="3" />
                    <RELAYPOSITION athleteid="36141" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="15. Deutsche Kurzbahnmeisterschaft der Masters" city="Essen" date="2025-11-30" qualificationtime="00:02:10.88" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="4">
              <ENTRIES>
                <ENTRY entrytime="00:02:31.99" eventid="1183" heatid="40143" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="36257" number="1" />
                    <RELAYPOSITION athleteid="36193" number="2" />
                    <RELAYPOSITION athleteid="36049" number="3" />
                    <RELAYPOSITION athleteid="36093" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="15. Deutsche Kurzbahnmeisterschaft der Masters" city="Essen" date="2025-11-30" qualificationtime="00:02:10.88" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="3332" nation="GER" region="12" clubid="39228" name="Dresdner SC 1898">
          <ATHLETES>
            <ATHLETE firstname="Bruno" lastname="Hutzler" birthdate="2010-01-01" gender="M" nation="GER" license="410638" athleteid="39588">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.78" eventid="1133" heatid="40074" lane="7">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:29.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.69" eventid="1237" heatid="40223" lane="5">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:15.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.04" eventid="1153" heatid="40107" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:02:47.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.52" eventid="1277" heatid="40298" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:01:04.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.36" eventid="1297" heatid="40338" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:31.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.30" eventid="1337" heatid="40398" lane="5">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:19.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.05" eventid="1217" heatid="40185" lane="5">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:34.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.03" eventid="1377" heatid="40467" lane="4">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:33.50" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Heidi" lastname="Hanel" birthdate="2012-01-01" gender="F" nation="GER" license="436913" athleteid="39606">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.88" eventid="1123" heatid="40046" lane="4">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:30.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.48" eventid="1267" heatid="40272" lane="6">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:10.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.97" eventid="1207" heatid="40163" lane="7">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:40.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.53" eventid="1367" heatid="40450" lane="1">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Kolkowski" birthdate="2012-01-01" gender="M" nation="GER" license="443040" athleteid="39655">
              <ENTRIES>
                <ENTRY entrytime="00:02:40.61" eventid="1197" heatid="40153" lane="4">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:02:40.61" />
                </ENTRY>
                <ENTRY entrytime="00:19:03.96" eventid="1113" heatid="40025" lane="8">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-14" qualificationtime="00:19:03.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.69" eventid="1277" heatid="40301" lane="1">
                  <MEETINFO name="DMSJ - Landesentscheid Sachsen" city="Dresden" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:01:02.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.67" eventid="1377" heatid="40470" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:31.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.57" eventid="1173" heatid="40138" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:24.66" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.62" eventid="1237" heatid="40228" lane="7">
                  <MEETINFO name="DMSJ - Landesentscheid Sachsen" city="Dresden" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:01:07.68" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.74" eventid="1397" heatid="40492" lane="1">
                  <MEETINFO name="DMSJ - Landesentscheid Sachsen" city="Dresden" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:01:07.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jasmin" lastname="Suha" birthdate="2013-01-01" gender="F" nation="GER" license="443682" athleteid="39800">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.30" eventid="1123" heatid="40028" lane="1">
                  <MEETINFO name="Stadtmeisterschaft Dresden" city="Dresden" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:36.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.98" eventid="1207" heatid="40159" lane="3" />
                <ENTRY entrytime="00:01:30.64" eventid="1227" heatid="40194" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:27.44" />
                </ENTRY>
                <ENTRY entrytime="00:03:17.86" eventid="1163" heatid="40113" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alexej" lastname="Chaplygin" birthdate="2012-01-01" gender="M" nation="GER" license="443662" athleteid="39290">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.73" eventid="1237" heatid="40222" lane="4">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:19.73" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.59" eventid="1357" heatid="40423" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:49.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.97" eventid="1377" heatid="40465" lane="3">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:00:36.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.42" eventid="1277" heatid="40295" lane="1">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:11.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.17" eventid="1217" heatid="40177" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:44.17" />
                </ENTRY>
                <ENTRY entrytime="00:06:03.64" eventid="1257" heatid="40247" lane="1">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:06:03.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.62" eventid="1337" heatid="40395" lane="8">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:01:32.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Greta" lastname="Bachmann" birthdate="2011-01-01" gender="F" nation="GER" license="424908" athleteid="39719">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.88" eventid="1123" heatid="40041" lane="1">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:31.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.61" eventid="1227" heatid="40204" lane="8">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:01:19.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Benno" lastname="Salfitzky" birthdate="2014-01-01" gender="M" nation="GER" license="448061" athleteid="39259">
              <ENTRIES>
                <ENTRY entrytime="00:02:30.07" eventid="1357" heatid="40427" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:27.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.87" eventid="1297" heatid="40337" lane="6">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:32.31" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.85" eventid="1257" heatid="40252" lane="2">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:05:15.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.43" eventid="1133" heatid="40075" lane="2">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:29.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.55" eventid="1277" heatid="40297" lane="4">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:05.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.53" eventid="1173" heatid="40138" lane="8">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:02:37.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Dunkel" birthdate="2010-01-01" gender="F" nation="GER" license="410626" athleteid="39764">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.87" eventid="1123" heatid="40032" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:33.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.33" eventid="1367" heatid="40452" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:35.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.57" eventid="1227" heatid="40204" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:19.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jonas" lastname="Dieckow" birthdate="1999-01-01" gender="M" nation="GER" license="202175" athleteid="39307">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.07" eventid="1133" heatid="40082" lane="3">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-31" qualificationtime="00:00:27.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.00" eventid="1173" heatid="40139" lane="7" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Niklas" lastname="Wiese" birthdate="2013-01-01" gender="M" nation="GER" license="445789" athleteid="39968">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.96" eventid="1277" heatid="40296" lane="2">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:09.96" />
                </ENTRY>
                <ENTRY entrytime="00:10:38.82" eventid="1093" heatid="40015" lane="8">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:10:38.82" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.82" eventid="1317" heatid="40370" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:40.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.28" eventid="1217" heatid="40179" lane="3">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:40.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.99" eventid="1237" heatid="40224" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:01:16.99" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.73" eventid="1173" heatid="40136" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:02:41.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.64" eventid="1377" heatid="40465" lane="5">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:36.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Janina" lastname="Pannasch" birthdate="2000-01-01" gender="F" nation="GER" license="240074" athleteid="39667">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.72" eventid="1367" heatid="40449" lane="3">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:00:36.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.18" eventid="1287" heatid="40322" lane="3">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:00:33.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Kruse" birthdate="2007-01-01" gender="M" nation="GER" license="364582" athleteid="39229">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.07" eventid="1133" heatid="40082" lane="5">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:27.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.14" eventid="1297" heatid="40341" lane="2">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:30.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.11" eventid="1217" heatid="40186" lane="3">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:34.11" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Ulbricht" birthdate="2013-01-01" gender="M" nation="GER" license="443686" athleteid="39674">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.19" eventid="1277" heatid="40289" lane="3">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:20.19" />
                </ENTRY>
                <ENTRY entrytime="00:05:40.98" eventid="1257" heatid="40248" lane="2">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:06:06.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.98" eventid="1337" heatid="40392" lane="3">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:41.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.29" eventid="1237" heatid="40216" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:29.15" />
                </ENTRY>
                <ENTRY entrytime="00:01:44.12" eventid="1397" heatid="40486" lane="3">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:43.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.46" eventid="1133" heatid="40062" lane="6">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:00:35.46" />
                </ENTRY>
                <ENTRY entrytime="00:03:19.66" eventid="1173" heatid="40128" lane="4">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:03:19.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Leuteritz" birthdate="2010-01-01" gender="F" nation="GER" license="436108" athleteid="39813">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.53" eventid="1367" heatid="40450" lane="7">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:36.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.67" eventid="1123" heatid="40043" lane="8">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:31.67" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.36" eventid="1267" heatid="40274" lane="6">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:09.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.45" eventid="1287" heatid="40317" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:35.45" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marie-Luise" lastname="Rießland" birthdate="2006-01-01" gender="F" nation="GER" license="357421" athleteid="39868">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.98" eventid="1123" heatid="40046" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:30.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.99" eventid="1367" heatid="40449" lane="2">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:37.50" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fabian" lastname="Schellhammer" birthdate="2015-01-01" gender="M" nation="GER" license="463209" athleteid="39944">
              <ENTRIES>
                <ENTRY entrytime="00:01:26.92" eventid="1277" heatid="40288" lane="8">
                  <MEETINFO name="Giraffenpokal" city="Chemnitz" course="LCM" approved="GER" date="2025-11-08" qualificationtime="00:01:26.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.00" eventid="1397" heatid="40486" lane="6" />
                <ENTRY entrytime="00:00:42.43" eventid="1377" heatid="40461" lane="6">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:41.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.97" eventid="1297" heatid="40332" lane="1">
                  <MEETINFO name="Giraffenpokal" city="Chemnitz" course="LCM" approved="GER" date="2025-11-08" qualificationtime="00:00:41.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.07" eventid="1133" heatid="40060" lane="4">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:37.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.24" eventid="1237" heatid="40215" lane="5">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:34.24" />
                </ENTRY>
                <ENTRY entrytime="00:03:19.00" eventid="1173" heatid="40129" lane="8">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:03:19.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Carlotta" lastname="Harnisch" birthdate="2014-01-01" gender="F" nation="GER" license="448039" athleteid="39844">
              <ENTRIES>
                <ENTRY entrytime="00:01:27.52" eventid="1227" heatid="40196" lane="7">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:27.52" />
                </ENTRY>
                <ENTRY entrytime="00:05:55.98" eventid="1247" heatid="40235" lane="7" />
                <ENTRY entrytime="00:00:34.60" eventid="1123" heatid="40031" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:34.60" />
                </ENTRY>
                <ENTRY entrytime="00:01:41.40" eventid="1327" heatid="40379" lane="7">
                  <MEETINFO name="12. Erich Kästner Schwimmfest" city="Dresden" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:41.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.13" eventid="1267" heatid="40265" lane="7">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:18.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.28" eventid="1367" heatid="40444" lane="2">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:39.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Theodor" lastname="Gruhl" birthdate="2013-01-01" gender="M" nation="GER" license="445434" athleteid="39334">
              <ENTRIES>
                <ENTRY entrytime="00:10:45.00" eventid="1093" heatid="40014" lane="6">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-26" qualificationtime="00:11:48.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.44" eventid="1297" heatid="40334" lane="4">
                  <MEETINFO name="33. Internationale Geraer Stadtmeisterschaften" city="Gera" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:00:35.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.07" eventid="1237" heatid="40220" lane="5">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:21.08" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.51" eventid="1257" heatid="40252" lane="6">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:15.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.88" eventid="1377" heatid="40464" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:36.82" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.34" eventid="1153" heatid="40105" lane="3">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:03:07.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.91" eventid="1337" heatid="40396" lane="8">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:28.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lydia" lastname="Brüll" birthdate="2015-01-01" gender="F" nation="GER" license="463215" athleteid="39483">
              <ENTRIES>
                <ENTRY entrytime="00:01:38.98" eventid="1227" heatid="40192" lane="7">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:38.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.21" eventid="1123" heatid="40027" lane="7">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:00:38.21" />
                </ENTRY>
                <ENTRY entrytime="00:06:15.98" eventid="1247" heatid="40234" lane="2" />
                <ENTRY entrytime="00:03:09.89" eventid="1347" heatid="40404" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:03:09.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.98" eventid="1327" heatid="40377" lane="5">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:01:59.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.70" eventid="1267" heatid="40262" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:23.70" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Charlotte" lastname="von Bonin" birthdate="2009-01-01" gender="F" nation="GER" license="393877" athleteid="39465">
              <ENTRIES>
                <ENTRY entrytime="00:01:22.35" eventid="1227" heatid="40200" lane="4">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:19.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.61" eventid="1367" heatid="40448" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:35.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.94" eventid="1287" heatid="40318" lane="6">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:34.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.99" eventid="1123" heatid="40040" lane="1">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:31.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.37" eventid="1163" heatid="40116" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:02:54.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fredo Matheo" lastname="Schiller" birthdate="2012-01-01" gender="M" nation="GER" license="436894" athleteid="39382">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.02" eventid="1297" heatid="40334" lane="7">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:36.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.58" eventid="1133" heatid="40065" lane="6">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:33.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.70" eventid="1277" heatid="40293" lane="8">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:15.70" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Cornelius" lastname="Schramm" birthdate="2004-01-01" gender="M" nation="GER" license="309882" athleteid="39391">
              <ENTRIES>
                <ENTRY entrytime="00:02:22.15" eventid="1173" heatid="40140" lane="3">
                  <MEETINFO name="39. Internationale DM Masters Lange Strecke" city="Wolfsburg" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:02:26.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.46" eventid="1133" heatid="40087" lane="2" />
                <ENTRY entrytime="00:02:20.93" eventid="1317" heatid="40375" lane="3">
                  <MEETINFO name="15. Deutsche Kurzbahnmeisterschaft der Masters" city="Essen" course="SCM" approved="GER" date="2025-11-28" qualificationtime="00:02:15.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.83" eventid="1237" heatid="40230" lane="4">
                  <MEETINFO name="15. Deutsche Kurzbahnmeisterschaft der Masters" city="Essen" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:01:00.97" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karl Hugo" lastname="Lages" birthdate="2015-01-01" gender="M" nation="GER" license="463216" athleteid="39429">
              <ENTRIES>
                <ENTRY entrytime="00:03:06.59" eventid="1357" heatid="40421" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:03:06.59" />
                </ENTRY>
                <ENTRY entrytime="00:03:49.14" eventid="1153" heatid="40101" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:03:49.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.75" eventid="1217" heatid="40175" lane="2">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:45.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.89" eventid="1237" heatid="40216" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:32.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:44.09" eventid="1337" heatid="40391" lane="5">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:44.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.71" eventid="1277" heatid="40288" lane="2">
                  <MEETINFO name="12. Erich Kästner Schwimmfest" city="Dresden" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:24.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Henrijette" lastname="Kobus" birthdate="2012-01-01" gender="F" nation="GER" license="439567" athleteid="39643">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.53" eventid="1367" heatid="40458" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:31.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.26" eventid="1123" heatid="40056" lane="6">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:00:28.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.63" eventid="1267" heatid="40283" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:01.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.11" eventid="1163" heatid="40126" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:22.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.18" eventid="1227" heatid="40212" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:06.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.83" eventid="1307" heatid="40360" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:33.83" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ferris" lastname="Winkler" birthdate="2008-01-01" gender="M" nation="GER" license="380816" athleteid="39952">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.20" eventid="1237" heatid="40228" lane="6">
                  <MEETINFO name="16. Internationales Nachwuchsschwimmfest" city="Cottbus" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:11.20" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.96" eventid="1217" heatid="40184" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:35.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.36" eventid="1277" heatid="40305" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:59.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.55" eventid="1133" heatid="40084" lane="3">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:25.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.04" eventid="1377" heatid="40472" lane="7">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:30.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.11" eventid="1297" heatid="40344" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:27.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.88" eventid="1397" heatid="40493" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:03.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Christian" lastname="Schubert" birthdate="2010-01-01" gender="M" nation="GER" license="412734" athleteid="39707">
              <ENTRIES>
                <ENTRY entrytime="00:04:09.34" eventid="1257" heatid="40260" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:04:09.34" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.95" eventid="1357" heatid="40438" lane="8">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:02:01.95" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.98" eventid="1317" heatid="40373" lane="5" />
                <ENTRY entrytime="00:02:21.37" eventid="1173" heatid="40140" lane="4" />
                <ENTRY entrytime="00:08:40.52" eventid="1093" heatid="40019" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:08:40.52" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Felix" lastname="Mehner" birthdate="2009-01-01" gender="M" nation="GER" license="395569" athleteid="39298">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.96" eventid="1237" heatid="40230" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:05.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.47" eventid="1397" heatid="40491" lane="7">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:01:11.47" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.28" eventid="1173" heatid="40139" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:31.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.70" eventid="1297" heatid="40342" lane="7">
                  <MEETINFO name="16. Internationales Nachwuchsschwimmfest" city="Cottbus" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:29.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.95" eventid="1133" heatid="40083" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:26.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.72" eventid="1277" heatid="40308" lane="1">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:57.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.48" eventid="1217" heatid="40183" lane="2">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:35.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.21" eventid="1377" heatid="40471" lane="4">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:30.52" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Friedrich" lastname="Deichmüller" birthdate="2015-01-01" gender="M" nation="GER" license="463211" athleteid="39878">
              <ENTRIES>
                <ENTRY entrytime="00:01:26.98" eventid="1277" heatid="40287" lane="3">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:01:30.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.98" eventid="1337" heatid="40391" lane="1">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:01:55.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.98" eventid="1377" heatid="40461" lane="5">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:41.96" />
                </ENTRY>
                <ENTRY entrytime="00:03:17.32" eventid="1173" heatid="40129" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:03:17.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.15" eventid="1237" heatid="40216" lane="2">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:01:32.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:49.98" eventid="1217" heatid="40174" lane="7">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:50.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Dörfer" birthdate="2009-01-01" gender="F" nation="GER" license="393881" athleteid="39342">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.95" eventid="1387" heatid="40481" lane="3">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:15.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.82" eventid="1287" heatid="40326" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:31.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.20" eventid="1227" heatid="40211" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:10.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.41" eventid="1123" heatid="40044" lane="7">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:30.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.16" eventid="1367" heatid="40458" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:30.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Florentine" lastname="Auerswald" birthdate="2011-01-01" gender="F" nation="GER" license="424902" athleteid="39818">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.99" eventid="1123" heatid="40030" lane="1">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:37.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.91" eventid="1207" heatid="40163" lane="3">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:41.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marie" lastname="Kruse" birthdate="2011-01-01" gender="F" nation="GER" license="424900" athleteid="39575">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.67" eventid="1367" heatid="40447" lane="4">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:37.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.10" eventid="1123" heatid="40045" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:31.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.10" eventid="1207" heatid="40162" lane="5">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:41.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.90" eventid="1267" heatid="40270" lane="5">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:01:11.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Erik" lastname="Dittmar" birthdate="2007-01-01" gender="M" nation="GER" license="364564" athleteid="39828">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.96" eventid="1297" heatid="40343" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:28.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.02" eventid="1277" heatid="40305" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:57.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.33" eventid="1217" heatid="40185" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.00" eventid="1377" heatid="40472" lane="2">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:29.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.26" eventid="1133" heatid="40082" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:26.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.89" eventid="1357" heatid="40432" lane="5">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:02:10.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.78" eventid="1173" heatid="40137" lane="4">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:02:37.78" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Levi" lastname="Martin" birthdate="2010-01-01" gender="M" nation="GER" license="424888" athleteid="39279">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.50" eventid="1277" heatid="40296" lane="6">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:09.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.59" eventid="1133" heatid="40072" lane="8">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:30.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.46" eventid="1217" heatid="40183" lane="6">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:36.46" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Klara" lastname="Beckmann" birthdate="2015-01-01" gender="F" nation="GER" license="463195" athleteid="39768">
              <ENTRIES>
                <ENTRY entrytime="00:03:27.65" eventid="1163" heatid="40112" lane="3">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:03:27.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:39.73" eventid="1227" heatid="40192" lane="1">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:39.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.98" eventid="1267" heatid="40261" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:30.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:47.78" eventid="1327" heatid="40378" lane="2">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:47.78" />
                </ENTRY>
                <ENTRY entrytime="00:06:15.98" eventid="1247" heatid="40234" lane="7" />
                <ENTRY entrytime="00:00:46.98" eventid="1367" heatid="40439" lane="5">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:44.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Rößler" birthdate="1997-01-01" gender="F" nation="GER" license="181670" athleteid="39357">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.72" eventid="1387" heatid="40479" lane="3">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:21.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.68" eventid="1347" heatid="40413" lane="6">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-31" qualificationtime="00:02:30.96" />
                </ENTRY>
                <ENTRY entrytime="00:19:44.82" eventid="1103" heatid="40021" lane="6">
                  <MEETINFO name="39. Internationale DM Masters Lange Strecke" city="Wolfsburg" course="LCM" approved="GER" date="2025-03-14" qualificationtime="00:21:42.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.36" eventid="1327" heatid="40385" lane="2">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:24.60" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.07" eventid="1267" heatid="40277" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:07.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Gähler" birthdate="2005-01-01" gender="M" nation="GER" license="349776" athleteid="39788">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.99" eventid="1133" heatid="40076" lane="2">
                  <MEETINFO name="28. Internationaler Sportbadpokal" city="Berlin" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:00:29.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.99" eventid="1377" heatid="40468" lane="8">
                  <MEETINFO name="28. Internationaler Sportbadpokal" city="Berlin" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:00:36.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Sachse" birthdate="2008-01-01" gender="M" nation="GER" license="380809" athleteid="39403">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.91" eventid="1297" heatid="40341" lane="3">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:29.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.94" eventid="1133" heatid="40083" lane="3">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:26.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.39" eventid="1337" heatid="40399" lane="2">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:16.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.51" eventid="1217" heatid="40186" lane="1">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:33.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.08" eventid="1377" heatid="40468" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:34.08" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.82" eventid="1397" heatid="40492" lane="2">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:06.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karl" lastname="Fritzsche" birthdate="2012-01-01" gender="M" nation="GER" license="445371" athleteid="39522">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.59" eventid="1237" heatid="40222" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:20.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.96" eventid="1337" heatid="40395" lane="2">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:29.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.80" eventid="1133" heatid="40067" lane="2">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:32.80" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Kirsten" birthdate="2014-01-01" gender="F" nation="GER" license="448042" athleteid="39533">
              <ENTRIES>
                <ENTRY entrytime="00:02:49.90" eventid="1163" heatid="40120" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:02:49.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.11" eventid="1347" heatid="40408" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:44.11" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.10" eventid="1307" heatid="40353" lane="2">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:54.82" />
                </ENTRY>
                <ENTRY entrytime="00:05:39.28" eventid="1247" heatid="40236" lane="3">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:05:39.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.23" eventid="1227" heatid="40203" lane="2">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:15.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.30" eventid="1123" heatid="40031" lane="5">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:33.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.79" eventid="1267" heatid="40269" lane="7">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:12.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Haufe" birthdate="2009-01-01" gender="M" nation="GER" license="410632" athleteid="39273">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.29" eventid="1133" heatid="40081" lane="5">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:27.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.27" eventid="1397" heatid="40492" lane="5">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:08.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.79" eventid="1297" heatid="40343" lane="5">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:28.79" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.62" eventid="1277" heatid="40302" lane="5">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:01:02.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.62" eventid="1237" heatid="40227" lane="7">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:12.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ella" lastname="Kirchner" birthdate="2015-01-01" gender="F" nation="GER" license="463200" athleteid="39912">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.86" eventid="1123" heatid="40036" lane="1">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:31.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.47" eventid="1163" heatid="40116" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:59.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.27" eventid="1267" heatid="40270" lane="7">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:09.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.43" eventid="1307" heatid="40352" lane="8">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:02:59.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.43" eventid="1227" heatid="40201" lane="4">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:21.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.22" eventid="1207" heatid="40160" lane="2">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:42.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.09" eventid="1367" heatid="40447" lane="1">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:36.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.15" eventid="1387" heatid="40477" lane="8">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:31.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Miriam" lastname="Junge" birthdate="2008-01-01" gender="F" nation="GER" license="390588" athleteid="39379">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.99" eventid="1123" heatid="40035" lane="5">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:32.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.57" eventid="1207" heatid="40166" lane="1">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:41.87" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Pepe Luis" lastname="Mattke" birthdate="2015-01-01" gender="M" nation="GER" license="463212" athleteid="39509">
              <ENTRIES>
                <ENTRY entrytime="00:03:05.80" eventid="1173" heatid="40130" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:03:05.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.07" eventid="1237" heatid="40219" lane="6">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:01:25.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.01" eventid="1277" heatid="40289" lane="5">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:01:20.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.90" eventid="1297" heatid="40333" lane="7">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:37.05" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.69" eventid="1133" heatid="40063" lane="6">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:34.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.32" eventid="1377" heatid="40464" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:38.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.46" eventid="1357" heatid="40423" lane="2">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:51.46" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ben" lastname="Gruner" birthdate="2009-01-01" gender="M" nation="GER" license="380717" athleteid="39497">
              <ENTRIES>
                <ENTRY entrytime="00:01:21.91" eventid="1337" heatid="40397" lane="4">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:18.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.10" eventid="1297" heatid="40340" lane="1">
                  <MEETINFO name="Stadtmeisterschaft Dresden" city="Dresden" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:31.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.12" eventid="1133" heatid="40076" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:28.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.00" eventid="1217" heatid="40184" lane="6">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:36.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alexandra" lastname="Kirberger" birthdate="2012-01-01" gender="F" nation="GER" license="436906" athleteid="39744">
              <ENTRIES>
                <ENTRY entrytime="00:05:46.09" eventid="1063" heatid="39996" lane="7">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-26" qualificationtime="00:05:46.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.64" eventid="1387" heatid="40484" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:09.53" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.27" eventid="1347" heatid="40417" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:18.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.89" eventid="1287" heatid="40328" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:30.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.81" eventid="1163" heatid="40124" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:30.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.82" eventid="1187" heatid="40149" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:29.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jonathan" lastname="Korn" birthdate="2006-01-01" gender="M" nation="GER" license="349797" athleteid="39517">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.05" eventid="1133" heatid="40082" lane="4">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:00:26.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.26" eventid="1297" heatid="40342" lane="4">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:00:28.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.50" eventid="1217" heatid="40187" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:33.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.93" eventid="1337" heatid="40399" lane="7">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:14.87" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Lieske" birthdate="2015-01-01" gender="M" nation="GER" license="463225" athleteid="39729">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.07" eventid="1133" heatid="40059" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:41.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.91" eventid="1377" heatid="40461" lane="8">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:45.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Annika Loreen" lastname="Zische" birthdate="2009-01-01" gender="F" nation="GER" license="393879" athleteid="39618">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.82" eventid="1327" heatid="40390" lane="4">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:12.93" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.10" eventid="1307" heatid="40361" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:26.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.45" eventid="1387" heatid="40485" lane="3">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:04.25" />
                </ENTRY>
                <ENTRY entrytime="00:05:19.83" eventid="1063" heatid="39997" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-26" qualificationtime="00:05:19.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.00" eventid="1207" heatid="40173" lane="5">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:33.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.42" eventid="1143" heatid="40099" lane="1">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:47.42" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Amelie" lastname="Ritter" birthdate="2003-01-01" gender="F" nation="GER" license="315370" athleteid="39386">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.07" eventid="1287" heatid="40328" lane="1">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-30" qualificationtime="00:00:31.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.63" eventid="1123" heatid="40055" lane="3">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-31" qualificationtime="00:00:29.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.40" eventid="1163" heatid="40122" lane="1" />
                <ENTRY entrytime="00:01:02.50" eventid="1267" heatid="40284" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anne-Felicia" lastname="Wagenknecht" birthdate="2009-01-01" gender="F" nation="GER" license="395546" athleteid="39451">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.15" eventid="1227" heatid="40203" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:17.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.54" eventid="1347" heatid="40410" lane="5">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:37.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.94" eventid="1267" heatid="40272" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:01:09.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.99" eventid="1123" heatid="40039" lane="4">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:31.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Cedric" lastname="Banek" birthdate="2013-01-01" gender="M" nation="GER" license="460089" athleteid="39663">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.75" eventid="1377" heatid="40462" lane="3">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:40.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.98" eventid="1337" heatid="40393" lane="5">
                  <MEETINFO name="BaWü &amp; Süddt Meisterschaften SMK" city="Stuttgart" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:01:34.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.85" eventid="1133" heatid="40064" lane="4">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.40" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leonie" lastname="Glasewald" birthdate="2005-01-01" gender="F" nation="GER" license="340499" athleteid="39686">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.08" eventid="1287" heatid="40328" lane="8">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-30" qualificationtime="00:00:31.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.34" eventid="1123" heatid="40053" lane="3">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-31" qualificationtime="00:00:29.39" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.88" eventid="1387" heatid="40483" lane="3">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:10.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.74" eventid="1367" heatid="40457" lane="4">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-06-01" qualificationtime="00:00:33.21" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.29" eventid="1227" heatid="40211" lane="8">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:09.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Pia" lastname="Müller" birthdate="2014-01-01" gender="F" nation="GER" license="448027" athleteid="39976">
              <ENTRIES>
                <ENTRY entrytime="00:02:43.98" eventid="1347" heatid="40408" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:43.98" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.29" eventid="1267" heatid="40274" lane="3">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:08.43" />
                </ENTRY>
                <ENTRY entrytime="00:03:04.59" eventid="1163" heatid="40115" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:03:04.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.80" eventid="1307" heatid="40352" lane="4">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:54.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.20" eventid="1207" heatid="40159" lane="7">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:43.68" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.12" eventid="1227" heatid="40199" lane="5">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:20.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.01" eventid="1123" heatid="40035" lane="3">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:31.45" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Kiss" birthdate="2011-01-01" gender="F" nation="GER" license="448034" athleteid="39348">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.57" eventid="1123" heatid="40037" lane="8">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:32.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.88" eventid="1287" heatid="40316" lane="4">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:00:35.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.98" eventid="1267" heatid="40270" lane="3">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:01:11.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.10" eventid="1367" heatid="40447" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:38.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Konstantin" lastname="Silex" birthdate="2008-01-01" gender="M" nation="GER" license="387209" athleteid="39317">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.76" eventid="1173" heatid="40142" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:06.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.08" eventid="1377" heatid="40474" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:27.80" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.47" eventid="1317" heatid="40376" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:15.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.35" eventid="1237" heatid="40232" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:59.26" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Peter" lastname="Dürrling" birthdate="2007-01-01" gender="M" nation="GER" license="380795" athleteid="39775">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.21" eventid="1297" heatid="40338" lane="4">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:31.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.24" eventid="1217" heatid="40185" lane="3">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.08" eventid="1337" heatid="40398" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:16.61" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.22" eventid="1153" heatid="40106" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:02:54.56" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Julian" lastname="Nietzold" birthdate="2007-01-01" gender="M" nation="GER" license="364589" athleteid="39580">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.99" eventid="1133" heatid="40076" lane="7">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:29.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.99" eventid="1377" heatid="40468" lane="1">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:34.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Erik" lastname="Beckmann" birthdate="2015-01-01" gender="M" nation="GER" license="463196" athleteid="39921">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" eventid="1297" heatid="40332" lane="6">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:39.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.50" eventid="1133" heatid="40061" lane="6">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:35.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.93" eventid="1237" heatid="40215" lane="7">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:35.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.24" eventid="1337" heatid="40392" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:43.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.71" eventid="1277" heatid="40288" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:22.71" />
                </ENTRY>
                <ENTRY entrytime="00:03:30.98" eventid="1173" heatid="40128" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:03:31.80" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Schwöd" birthdate="2006-01-01" gender="F" nation="GER" license="370572" athleteid="39322">
              <ENTRIES>
                <ENTRY entrytime="00:03:06.00" eventid="1143" heatid="40095" lane="5">
                  <MEETINFO name="DMS-Austragung 24/25 Bezirksliga - Oberpfalz" city="Weiden" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:02:59.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.00" eventid="1287" heatid="40323" lane="6">
                  <MEETINFO name="22. Internationales Landauer Dreikönigsschwimmen" city="Landau/Isar" course="SCM" approved="GER" date="2025-01-06" qualificationtime="00:00:32.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.90" eventid="1327" heatid="40387" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:21.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.77" eventid="1207" heatid="40169" lane="2">
                  <MEETINFO name="11. Wackersdorfer Panoramabadschwimmfest" city="Wackersdorf" course="SCM" approved="GER" date="2025-07-12" qualificationtime="00:00:37.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.29" eventid="1387" heatid="40482" lane="7">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:11.66" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.00" eventid="1227" heatid="40203" lane="3">
                  <MEETINFO name="25. Internationales Landauer Sprinter-Treffen" city="Landau/Isar" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:13.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mathilde" lastname="Brendler" birthdate="2008-01-01" gender="F" nation="GER" license="380792" athleteid="39363">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.27" eventid="1287" heatid="40320" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:34.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.30" eventid="1367" heatid="40450" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:36.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.26" eventid="1123" heatid="40044" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:31.26" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Stange" birthdate="2012-01-01" gender="F" nation="GER" license="436920" athleteid="39751">
              <ENTRIES>
                <ENTRY entrytime="00:01:16.98" eventid="1267" heatid="40265" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:22.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.98" eventid="1207" heatid="40160" lane="6">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:49.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.98" eventid="1123" heatid="40028" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:37.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.98" eventid="1327" heatid="40380" lane="7">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:43.67" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.73" eventid="1227" heatid="40194" lane="5">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:30.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.34" eventid="1367" heatid="40442" lane="3">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:40.34" />
                </ENTRY>
                <ENTRY entrytime="00:03:15.98" eventid="1163" heatid="40113" lane="3">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:03:23.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Artem" lastname="Lukasevych" birthdate="2010-01-01" gender="M" nation="GER" license="456870" athleteid="39233">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.20" eventid="1217" heatid="40182" lane="3">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:36.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.64" eventid="1397" heatid="40490" lane="4">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:01:14.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.06" eventid="1277" heatid="40302" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:03.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.81" eventid="1297" heatid="40338" lane="1">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:31.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.40" eventid="1377" heatid="40471" lane="8">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:31.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.88" eventid="1237" heatid="40228" lane="8">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:01:11.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.55" eventid="1133" heatid="40077" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:28.23" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Bastian" lastname="Höhne" birthdate="2006-01-01" gender="M" nation="GER" license="349790" athleteid="39625">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.82" eventid="1133" heatid="40076" lane="5">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:28.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.50" eventid="1237" heatid="40226" lane="1">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:12.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.85" eventid="1377" heatid="40470" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.11" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hannes" lastname="Winkler" birthdate="2011-01-01" gender="M" nation="GER" license="424910" athleteid="39597">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.99" eventid="1133" heatid="40069" lane="7">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:33.09" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Elena" lastname="Packenius" birthdate="2009-01-01" gender="F" nation="GER" license="396078" athleteid="39502">
              <ENTRIES>
                <ENTRY entrytime="00:02:50.51" eventid="1163" heatid="40119" lane="2">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:02:50.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.30" eventid="1287" heatid="40322" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:32.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.12" eventid="1123" heatid="40039" lane="1">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.98" eventid="1227" heatid="40206" lane="7">
                  <MEETINFO name="16. Internationales Nachwuchsschwimmfest" city="Cottbus" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:16.98" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.81" eventid="1387" heatid="40479" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:01:19.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.12" eventid="1367" heatid="40453" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Merle" lastname="Stange" birthdate="2015-01-01" gender="F" nation="GER" license="463204" athleteid="39890">
              <ENTRIES>
                <ENTRY entrytime="00:05:50.98" eventid="1143" heatid="40090" lane="8" />
                <ENTRY entrytime="00:01:26.98" eventid="1267" heatid="40261" lane="3">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:49.79" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.98" eventid="1227" heatid="40191" lane="4">
                  <MEETINFO name="12. Erich Kästner Schwimmfest" city="Dresden" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:44.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.61" eventid="1367" heatid="40440" lane="1">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:00:46.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.98" eventid="1327" heatid="40377" lane="4">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:02:01.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.98" eventid="1123" heatid="40026" lane="1">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:47.23" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Giesecke" birthdate="2009-01-01" gender="M" nation="GER" license="410628" athleteid="39423">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.47" eventid="1237" heatid="40226" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:11.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.11" eventid="1133" heatid="40079" lane="2">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:27.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.59" eventid="1277" heatid="40301" lane="7">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:01.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.21" eventid="1297" heatid="40341" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:29.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.45" eventid="1377" heatid="40470" lane="8">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Charlotte" lastname="Streiber" birthdate="2009-01-01" gender="F" nation="GER" license="398189" athleteid="39253">
              <ENTRIES>
                <ENTRY entrytime="00:02:29.17" eventid="1347" heatid="40414" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:02:39.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.07" eventid="1123" heatid="40045" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:30.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.48" eventid="1267" heatid="40274" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:01:09.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.49" eventid="1287" heatid="40319" lane="2">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:33.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.50" eventid="1227" heatid="40202" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:18.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Quentin" lastname="Schramm" birthdate="2007-01-01" gender="M" nation="GER" license="391015" athleteid="39546">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.07" eventid="1337" heatid="40399" lane="5">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:14.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.88" eventid="1133" heatid="40083" lane="4">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:26.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.01" eventid="1397" heatid="40493" lane="2">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:06.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.89" eventid="1217" heatid="40186" lane="4">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:33.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.10" eventid="1377" heatid="40468" lane="5">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:32.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.16" eventid="1297" heatid="40344" lane="7">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:28.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Uebel" birthdate="2015-01-01" gender="F" nation="GER" license="463205" athleteid="39241">
              <ENTRIES>
                <ENTRY entrytime="00:01:33.80" eventid="1227" heatid="40193" lane="5">
                  <MEETINFO name="12. Erich Kästner Schwimmfest" city="Dresden" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:33.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:42.42" eventid="1327" heatid="40379" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:42.42" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.74" eventid="1347" heatid="40405" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:03:01.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.37" eventid="1267" heatid="40264" lane="3">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:19.37" />
                </ENTRY>
                <ENTRY entrytime="00:03:40.08" eventid="1143" heatid="40090" lane="6">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:03:40.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.12" eventid="1123" heatid="40028" lane="2">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:34.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Felix" lastname="Kluge" birthdate="2014-01-01" gender="M" nation="GER" license="449664" athleteid="39905">
              <ENTRIES>
                <ENTRY entrytime="00:03:41.87" eventid="1153" heatid="40102" lane="1" />
                <ENTRY entrytime="00:01:18.01" eventid="1277" heatid="40291" lane="8">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:16.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.75" eventid="1297" heatid="40333" lane="3">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:00:36.75" />
                </ENTRY>
                <ENTRY entrytime="00:05:55.98" eventid="1257" heatid="40247" lane="2">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:06:06.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:41.92" eventid="1337" heatid="40392" lane="2">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:40.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.92" eventid="1237" heatid="40220" lane="8">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:23.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Göhre" birthdate="2014-01-01" gender="F" nation="GER" license="448209" athleteid="39821">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.84" eventid="1123" heatid="40033" lane="8">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:33.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.18" eventid="1227" heatid="40193" lane="2">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:35.18" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.98" eventid="1347" heatid="40404" lane="4">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:03:18.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.98" eventid="1327" heatid="40378" lane="3">
                  <MEETINFO name="12. Erich Kästner Schwimmfest" city="Dresden" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:02:05.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.39" eventid="1267" heatid="40263" lane="6">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:20.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.98" eventid="1207" heatid="40158" lane="8">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:52.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mateo" lastname="Blasius" birthdate="2010-01-01" gender="M" nation="GER" license="410623" athleteid="39561">
              <ENTRIES>
                <ENTRY entrytime="00:01:16.63" eventid="1237" heatid="40224" lane="5">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:01:16.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.87" eventid="1133" heatid="40073" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:28.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.82" eventid="1377" heatid="40469" lane="2">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:33.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.36" eventid="1297" heatid="40337" lane="1">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.64" eventid="1277" heatid="40297" lane="1">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:01:06.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Helen Ronja" lastname="Hein" birthdate="2014-01-01" gender="F" nation="GER" license="448835" athleteid="39936">
              <ENTRIES>
                <ENTRY entrytime="00:01:22.20" eventid="1227" heatid="40201" lane="7">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:01:22.20" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.27" eventid="1163" heatid="40118" lane="7">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:02:54.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.16" eventid="1347" heatid="40409" lane="7">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:02:41.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.55" eventid="1307" heatid="40353" lane="1">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:56.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.02" eventid="1367" heatid="40444" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:37.12" />
                </ENTRY>
                <ENTRY entrytime="00:11:40.00" eventid="1083" heatid="40004" lane="6">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:12:50.56" />
                </ENTRY>
                <ENTRY entrytime="00:05:36.15" eventid="1247" heatid="40237" lane="2">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:05:36.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jasmin" lastname="Zesewitz" birthdate="2006-01-01" gender="F" nation="GER" license="354302" athleteid="39471">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.66" eventid="1207" heatid="40171" lane="2">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:39.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.37" eventid="1347" heatid="40413" lane="5">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:02:33.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.26" eventid="1267" heatid="40278" lane="3" />
                <ENTRY entrytime="00:01:26.88" eventid="1327" heatid="40386" lane="1">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:30.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.18" eventid="1123" heatid="40049" lane="2">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:00:31.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Robin" lastname="Franke" birthdate="2015-01-01" gender="M" nation="GER" license="463214" athleteid="39541">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.68" eventid="1133" heatid="40061" lane="2">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:35.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:49.34" eventid="1217" heatid="40174" lane="3">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:49.34" />
                </ENTRY>
                <ENTRY entrytime="00:03:29.88" eventid="1173" heatid="40128" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:03:29.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:38.50" eventid="1237" heatid="40215" lane="8">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:01:38.50" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Franziska" lastname="Kirberger" birthdate="2015-01-01" gender="F" nation="GER" license="463223" athleteid="39791">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.34" eventid="1367" heatid="40441" lane="5">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:38.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.89" eventid="1123" heatid="40028" lane="3">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:33.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.52" eventid="1287" heatid="40313" lane="7">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:36.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.40" eventid="1387" heatid="40477" lane="6">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:29.40" />
                </ENTRY>
                <ENTRY entrytime="00:03:08.88" eventid="1163" heatid="40114" lane="7">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:03:08.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.33" eventid="1207" heatid="40158" lane="7">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:44.00" />
                </ENTRY>
                <ENTRY entrytime="00:03:06.06" eventid="1307" heatid="40350" lane="2">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:03:06.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.19" eventid="1227" heatid="40193" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:33.19" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Yanic" lastname="Paris" birthdate="2013-01-01" gender="M" nation="GER" license="448044" athleteid="39836">
              <ENTRIES>
                <ENTRY entrytime="00:03:08.84" eventid="1173" heatid="40130" lane="1">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:03:08.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.46" eventid="1297" heatid="40333" lane="6">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:37.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.98" eventid="1217" heatid="40177" lane="8">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:49.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.02" eventid="1277" heatid="40290" lane="4">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:18.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.48" eventid="1237" heatid="40217" lane="1">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:30.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.20" eventid="1377" heatid="40463" lane="8">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:40.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.98" eventid="1337" heatid="40392" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:45.68" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alissa" lastname="Ponomarenko" birthdate="2013-01-01" gender="F" nation="GER" license="443680" athleteid="39410">
              <ENTRIES>
                <ENTRY entrytime="00:03:20.98" eventid="1163" heatid="40113" lane="1" />
                <ENTRY entrytime="00:00:36.12" eventid="1123" heatid="40028" lane="7">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:36.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.98" eventid="1327" heatid="40379" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:58.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.86" eventid="1227" heatid="40194" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:29.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.98" eventid="1267" heatid="40263" lane="1">
                  <MEETINFO name="12. Erich Kästner Schwimmfest" city="Dresden" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:21.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.98" eventid="1287" heatid="40312" lane="5">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:42.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.98" eventid="1367" heatid="40441" lane="2">
                  <MEETINFO name="Stadtmeisterschaft Dresden" city="Dresden" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:43.44" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Felix" lastname="Müller" birthdate="2014-01-01" gender="M" nation="GER" license="447956" athleteid="39436">
              <ENTRIES>
                <ENTRY entrytime="00:01:24.92" eventid="1237" heatid="40219" lane="3">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:17.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.72" eventid="1133" heatid="40074" lane="6">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:29.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.77" eventid="1297" heatid="40336" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:33.76" />
                </ENTRY>
                <ENTRY entrytime="00:06:00.45" eventid="1073" heatid="39999" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:06:00.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.98" eventid="1397" heatid="40490" lane="5">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:01:14.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.28" eventid="1357" heatid="40429" lane="5">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:24.28" />
                </ENTRY>
                <ENTRY entrytime="00:05:24.06" eventid="1257" heatid="40250" lane="5">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:24.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Granzow" birthdate="2014-01-01" gender="M" nation="GER" license="448232" athleteid="39732">
              <ENTRIES>
                <ENTRY entrytime="00:01:34.99" eventid="1237" heatid="40215" lane="6">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:34.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.98" eventid="1217" heatid="40175" lane="1">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:52.57" />
                </ENTRY>
                <ENTRY entrytime="00:03:25.98" eventid="1173" heatid="40128" lane="2" />
                <ENTRY entrytime="00:00:36.94" eventid="1133" heatid="40061" lane="8">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:36.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Lange" birthdate="2013-01-01" gender="M" nation="GER" license="443672" athleteid="39928">
              <ENTRIES>
                <ENTRY entrytime="00:01:18.48" eventid="1397" heatid="40490" lane="8">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:01:18.48" />
                </ENTRY>
                <ENTRY entrytime="00:05:01.88" eventid="1257" heatid="40254" lane="4">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:01.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.30" eventid="1173" heatid="40137" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:35.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.73" eventid="1237" heatid="40225" lane="2">
                  <MEETINFO name="DMSJ - Landesentscheid Sachsen" city="Dresden" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:01:12.12" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.90" eventid="1357" heatid="40429" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:21.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.49" eventid="1133" heatid="40075" lane="1">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:29.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.25" eventid="1297" heatid="40338" lane="5">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:00:32.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Grischa" lastname="Ulbrich" birthdate="2011-01-01" gender="M" nation="GER" license="449835" athleteid="39698">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.99" eventid="1133" heatid="40069" lane="8">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.50" eventid="1237" heatid="40219" lane="1">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:22.40" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Schramm" birthdate="2012-01-01" gender="F" nation="GER" license="436911" athleteid="39418">
              <ENTRIES>
                <ENTRY entrytime="00:01:16.99" eventid="1267" heatid="40265" lane="5">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:17.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.95" eventid="1367" heatid="40445" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:38.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.40" eventid="1287" heatid="40316" lane="8">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:00:36.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.92" eventid="1123" heatid="40032" lane="5">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:33.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mattea" lastname="Schubert" birthdate="2007-01-01" gender="F" nation="GER" license="380811" athleteid="39288">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.59" eventid="1123" heatid="40058" lane="3">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:00:26.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Aurel" lastname="Wüstenhagen" birthdate="2009-01-01" gender="M" nation="GER" license="395576" athleteid="39329">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.74" eventid="1197" heatid="40156" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:07.64" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.75" eventid="1357" heatid="40436" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:01.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.18" eventid="1397" heatid="40496" lane="4">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:59.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.27" eventid="1317" heatid="40374" lane="6">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:23.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anna Lena" lastname="Gutjahr" birthdate="2014-01-01" gender="F" nation="GER" license="448021" athleteid="39310">
              <ENTRIES>
                <ENTRY entrytime="00:01:23.11" eventid="1227" heatid="40199" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:18.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.78" eventid="1123" heatid="40042" lane="1">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:31.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.32" eventid="1163" heatid="40118" lane="1">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:02:54.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.15" eventid="1367" heatid="40451" lane="8">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:00:35.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.00" eventid="1267" heatid="40273" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:09.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.01" eventid="1287" heatid="40323" lane="1">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:33.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nora" lastname="Fischer" birthdate="2015-01-01" gender="F" nation="GER" license="465835" athleteid="39851">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.71" eventid="1267" heatid="40268" lane="2">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:13.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.37" eventid="1123" heatid="40029" lane="3">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:32.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.13" eventid="1307" heatid="40353" lane="7">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:51.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.36" eventid="1387" heatid="40477" lane="3">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:29.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.61" eventid="1207" heatid="40161" lane="8">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:42.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.74" eventid="1227" heatid="40197" lane="8">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:25.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.87" eventid="1367" heatid="40443" lane="2">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:38.71" />
                </ENTRY>
                <ENTRY entrytime="00:03:06.99" eventid="1163" heatid="40114" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:03:06.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fynn Mario" lastname="Drzymala" birthdate="2008-01-01" gender="M" nation="GER" license="380796" athleteid="39713">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.77" eventid="1297" heatid="40346" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:26.17" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.99" eventid="1397" heatid="40495" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:58.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.10" eventid="1133" heatid="40085" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:25.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.24" eventid="1317" heatid="40375" lane="6" />
                <ENTRY entrytime="00:02:19.41" eventid="1197" heatid="40155" lane="5">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-25" qualificationtime="00:02:19.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mila" lastname="Mauermann" birthdate="2011-01-01" gender="F" nation="GER" license="424568" athleteid="39526">
              <ENTRIES>
                <ENTRY entrytime="00:04:37.10" eventid="1247" heatid="40245" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:04:37.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.37" eventid="1267" heatid="40285" lane="6">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:01:01.37" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.35" eventid="1387" heatid="40485" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:06.10" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.67" eventid="1347" heatid="40419" lane="4">
                  <MEETINFO name="Int. BAUAkademie ATUS Graz Trophy" city="Graz" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:02:13.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.63" eventid="1123" heatid="40055" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:28.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.19" eventid="1187" heatid="40150" lane="3">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:02:30.19" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Moritz" lastname="Haase" birthdate="2001-01-01" gender="M" nation="GER" license="261605" athleteid="39885">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.01" eventid="1237" heatid="40231" lane="1" />
                <ENTRY entrytime="00:00:54.02" eventid="1277" heatid="40311" lane="7" />
                <ENTRY entrytime="00:00:27.89" eventid="1377" heatid="40474" lane="6" />
                <ENTRY entrytime="00:00:24.88" eventid="1133" heatid="40088" lane="7" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Endrik" lastname="Böhme" birthdate="2015-01-01" gender="M" nation="GER" license="463193" athleteid="39599">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.98" eventid="1357" heatid="40421" lane="3" />
                <ENTRY entrytime="00:03:50.98" eventid="1153" heatid="40101" lane="5" />
                <ENTRY entrytime="00:01:50.98" eventid="1337" heatid="40391" lane="8">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:01:57.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:49.98" eventid="1217" heatid="40174" lane="2">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:52.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.98" eventid="1237" heatid="40214" lane="4">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:52.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.98" eventid="1277" heatid="40287" lane="4">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:52.49" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Timon" lastname="Böhme" birthdate="2012-01-01" gender="M" nation="GER" license="436922" athleteid="39367">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.85" eventid="1297" heatid="40337" lane="5">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:32.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.12" eventid="1277" heatid="40300" lane="5">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:04.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.64" eventid="1133" heatid="40077" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:28.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Martin" birthdate="2007-01-01" gender="M" nation="GER" license="364583" athleteid="39682">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.22" eventid="1377" heatid="40471" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:32.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.21" eventid="1133" heatid="40082" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:27.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.06" eventid="1297" heatid="40340" lane="7">
                  <MEETINFO name="28. Internationaler Sportbadpokal" city="Berlin" course="LCM" approved="GER" date="2025-06-08" qualificationtime="00:00:31.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Ritschel" birthdate="2007-01-01" gender="F" nation="GER" license="364594" athleteid="39960">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.60" eventid="1267" heatid="40280" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:04.37" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.74" eventid="1227" heatid="40202" lane="3">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:16.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.57" eventid="1123" heatid="40052" lane="6">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:29.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.26" eventid="1367" heatid="40453" lane="7">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.47" eventid="1207" heatid="40167" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:38.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.77" eventid="1387" heatid="40483" lane="4">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:01:11.77" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.44" eventid="1287" heatid="40327" lane="1">
                  <MEETINFO name="Sparkassen-Cup" city="Erlangen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:31.44" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mika-Frederik" lastname="Martin" birthdate="2012-01-01" gender="M" nation="GER" license="436899" athleteid="39371">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.18" eventid="1133" heatid="40085" lane="6">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:25.67" />
                </ENTRY>
                <ENTRY entrytime="00:04:23.64" eventid="1257" heatid="40259" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:04:23.64" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.09" eventid="1197" heatid="40155" lane="4">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:02:19.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.25" eventid="1357" heatid="40437" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:02:04.25" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.15" eventid="1397" heatid="40495" lane="3">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:00.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.10" eventid="1317" heatid="40374" lane="1">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:02:24.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.43" eventid="1277" heatid="40310" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:55.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Oliver" lastname="Manz" birthdate="1996-01-01" gender="M" nation="GER" license="181641" athleteid="39396">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.09" eventid="1377" heatid="40470" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:33.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jolien" lastname="Barthel-Krauße" birthdate="2014-01-01" gender="F" nation="GER" license="463382" athleteid="39490">
              <ENTRIES>
                <ENTRY entrytime="00:03:19.51" eventid="1163" heatid="40113" lane="7">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:03:19.51" />
                </ENTRY>
                <ENTRY entrytime="00:05:55.98" eventid="1247" heatid="40235" lane="1">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:06:44.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.26" eventid="1267" heatid="40262" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:23.26" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.98" eventid="1347" heatid="40405" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:03:07.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.98" eventid="1327" heatid="40378" lane="5">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:01:52.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.89" eventid="1227" heatid="40194" lane="1">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:32.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Henrik" lastname="Litta" birthdate="2015-01-01" gender="M" nation="GER" license="463806" athleteid="39456">
              <ENTRIES>
                <ENTRY entrytime="00:03:11.92" eventid="1173" heatid="40130" lane="8">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:03:11.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.55" eventid="1237" heatid="40218" lane="8">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:28.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.49" eventid="1277" heatid="40291" lane="5">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:16.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.22" eventid="1217" heatid="40176" lane="5">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:42.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.47" eventid="1377" heatid="40462" lane="5">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:40.26" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.30" eventid="1317" heatid="40364" lane="5">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:03:03.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.09" eventid="1337" heatid="40393" lane="3">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:32.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.01" eventid="1133" heatid="40061" lane="4">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:34.34" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Konstantin" lastname="Labuschke" birthdate="2014-01-01" gender="M" nation="GER" license="451949" athleteid="39860">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.03" eventid="1377" heatid="40461" lane="3">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:41.19" />
                </ENTRY>
                <ENTRY entrytime="00:03:41.87" eventid="1153" heatid="40102" lane="7" />
                <ENTRY entrytime="00:00:34.95" eventid="1133" heatid="40063" lane="2">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:34.90" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.98" eventid="1297" heatid="40331" lane="4">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:41.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.93" eventid="1277" heatid="40291" lane="6">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:16.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.20" eventid="1237" heatid="40216" lane="8">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:30.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.98" eventid="1337" heatid="40392" lane="8">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:43.78" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Scheffler" birthdate="2006-01-01" gender="F" nation="GER" license="353810" athleteid="39583">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.45" eventid="1123" heatid="40048" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:29.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.06" eventid="1367" heatid="40455" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:34.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.02" eventid="1207" heatid="40170" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:38.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.22" eventid="1287" heatid="40320" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:32.22" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alexandra" lastname="Schwendler" birthdate="2013-01-01" gender="F" nation="GER" license="449958" athleteid="39611">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.05" eventid="1367" heatid="40449" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:35.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.89" eventid="1227" heatid="40201" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:17.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.25" eventid="1123" heatid="40038" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:31.50" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.40" eventid="1347" heatid="40411" lane="5">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:35.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.05" eventid="1163" heatid="40118" lane="2">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:54.05" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.07" eventid="1287" heatid="40317" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:34.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Göde" birthdate="2008-01-01" gender="F" nation="GER" license="391855" athleteid="39692">
              <ENTRIES>
                <ENTRY entrytime="00:02:35.01" eventid="1307" heatid="40359" lane="4" />
                <ENTRY entrytime="00:01:04.58" eventid="1387" heatid="40485" lane="5">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:01:04.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.56" eventid="1123" heatid="40057" lane="3">
                  <MEETINFO name="Int. BAUAkademie ATUS Graz Trophy" city="Graz" course="LCM" approved="GER" date="2025-04-03" qualificationtime="00:00:27.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.41" eventid="1227" heatid="40212" lane="5">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:01:09.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.07" eventid="1267" heatid="40286" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:59.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hannah Victoria" lastname="Bürger" birthdate="2011-01-01" gender="F" nation="GER" license="424897" athleteid="39266">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.49" eventid="1367" heatid="40459" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:29.77" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.25" eventid="1123" heatid="40056" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.81" eventid="1163" heatid="40127" lane="4">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:02:21.81" />
                </ENTRY>
                <ENTRY entrytime="00:05:17.45" eventid="1063" heatid="39997" lane="7">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:05:17.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.21" eventid="1227" heatid="40213" lane="4">
                  <MEETINFO name="DMSJ - Landesentscheid Sachsen" city="Dresden" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:01:04.21" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.92" eventid="1307" heatid="40361" lane="3">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:24.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Frederike" lastname="Korn" birthdate="2010-01-01" gender="F" nation="GER" license="410641" athleteid="39759">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.13" eventid="1287" heatid="40316" lane="7">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:00:36.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.18" eventid="1123" heatid="40038" lane="4">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:32.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Adrian Leandro" lastname="Zische" birthdate="2008-01-01" gender="M" nation="GER" license="380817" athleteid="39248">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.13" eventid="1217" heatid="40189" lane="7">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:30.80" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.11" eventid="1153" heatid="40111" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:29.94" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.81" eventid="1357" heatid="40437" lane="2">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:02:04.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.79" eventid="1337" heatid="40402" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:06.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Matti" lastname="Ritschel" birthdate="2011-01-01" gender="M" nation="GER" license="424889" athleteid="39762">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.99" eventid="1133" heatid="40069" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:34.42" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maya" lastname="Tobehn" birthdate="2002-01-01" gender="F" nation="GER" license="292500" athleteid="39398">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.68" eventid="1267" heatid="40286" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:55.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.21" eventid="1287" heatid="40329" lane="4">
                  <MEETINFO name="Offene Finnische Meisterschaft" city="Helsinki" course="LCM" approved="GER" date="2025-06-26" qualificationtime="00:00:27.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.91" eventid="1123" heatid="40058" lane="4">
                  <MEETINFO name="Offene Finnische Meisterschaft" city="Helsinki" course="LCM" approved="GER" date="2025-06-27" qualificationtime="00:00:25.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.53" eventid="1347" heatid="40420" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:58.40" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Liepke" birthdate="2010-01-01" gender="M" nation="GER" license="397757" athleteid="39629">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.96" eventid="1297" heatid="40340" lane="3" />
                <ENTRY entrytime="00:02:13.85" eventid="1173" heatid="40142" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:09.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.67" eventid="1217" heatid="40188" lane="3">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:31.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.61" eventid="1133" heatid="40087" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:25.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.45" eventid="1237" heatid="40231" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:00.82" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.12" eventid="1357" heatid="40435" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:01.49" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.54" eventid="1317" heatid="40375" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:14.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leni" lastname="von Bonin" birthdate="2007-01-01" gender="F" nation="GER" license="364604" athleteid="39722">
              <ENTRIES>
                <ENTRY entrytime="00:08:45.31" eventid="1083" heatid="40011" lane="4">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:08:45.31" />
                </ENTRY>
                <ENTRY entrytime="00:04:09.57" eventid="1247" heatid="40245" lane="4">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:04:09.57" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="1227" heatid="40191" lane="3" />
                <ENTRY entrytime="00:02:26.62" eventid="1163" heatid="40127" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:18.61" />
                </ENTRY>
                <ENTRY entrytime="00:04:45.88" eventid="1063" heatid="39997" lane="4">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:04:40.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.02" eventid="1143" heatid="40099" lane="7" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Thorben" lastname="Salfitzky" birthdate="2010-01-01" gender="M" nation="GER" license="410651" athleteid="39871">
              <ENTRIES>
                <ENTRY entrytime="00:04:16.06" eventid="1257" heatid="40260" lane="8">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:04:16.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.50" eventid="1357" heatid="40437" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:00.25" />
                </ENTRY>
                <ENTRY entrytime="00:08:53.07" eventid="1093" heatid="40019" lane="1">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:08:53.07" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.24" eventid="1173" heatid="40141" lane="7">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:02:20.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.63" eventid="1277" heatid="40309" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:55.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.16" eventid="1317" heatid="40372" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nico" lastname="Koark" birthdate="2012-01-01" gender="M" nation="GER" license="436909" athleteid="39353">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.27" eventid="1133" heatid="40066" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:33.27" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.30" eventid="1237" heatid="40217" lane="7">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:30.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.99" eventid="1277" heatid="40292" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:16.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jakob" lastname="Schlott" birthdate="2009-01-01" gender="M" nation="GER" license="395539" athleteid="39477">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.74" eventid="1237" heatid="40228" lane="1">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:09.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.74" eventid="1133" heatid="40074" lane="2">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:29.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.68" eventid="1297" heatid="40339" lane="3">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:30.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.61" eventid="1377" heatid="40470" lane="5">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.96" eventid="1173" heatid="40136" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Hanke" birthdate="2010-01-01" gender="M" nation="GER" license="444305" athleteid="39650">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.00" eventid="1377" heatid="40466" lane="3">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:33.90" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.34" eventid="1297" heatid="40338" lane="3">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:32.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.88" eventid="1133" heatid="40073" lane="2">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:29.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.27" eventid="1217" heatid="40181" lane="6">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:38.24" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maike" lastname="Winkler" birthdate="2011-01-01" gender="F" nation="GER" license="424911" athleteid="39737">
              <ENTRIES>
                <ENTRY entrytime="00:02:28.81" eventid="1307" heatid="40361" lane="1">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:02:28.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.33" eventid="1387" heatid="40485" lane="6">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:01:06.33" />
                </ENTRY>
                <ENTRY entrytime="00:04:46.48" eventid="1247" heatid="40244" lane="4">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:04:46.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.21" eventid="1287" heatid="40329" lane="2">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:00:29.21" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.69" eventid="1267" heatid="40285" lane="5">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:01:00.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.05" eventid="1123" heatid="40058" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:26.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ria Johanna" lastname="Plietker" birthdate="2014-01-01" gender="F" nation="GER" license="448836" athleteid="39567">
              <ENTRIES>
                <ENTRY entrytime="00:01:21.28" eventid="1267" heatid="40263" lane="8">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:21.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.37" eventid="1227" heatid="40194" lane="2">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:32.37" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.78" eventid="1123" heatid="40028" lane="5">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:35.29" />
                </ENTRY>
                <ENTRY entrytime="00:03:39.71" eventid="1143" heatid="40090" lane="3">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:03:39.71" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.31" eventid="1327" heatid="40380" lane="5">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:01:35.31" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.98" eventid="1347" heatid="40404" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:03:08.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.37" eventid="1207" heatid="40161" lane="7">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:43.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marec Moritz" lastname="Pöschmann" birthdate="2009-01-01" gender="M" nation="GER" license="415182" athleteid="39637">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.49" eventid="1357" heatid="40438" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:55.94" />
                </ENTRY>
                <ENTRY entrytime="00:04:10.22" eventid="1257" heatid="40260" lane="2">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:04:10.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.77" eventid="1173" heatid="40141" lane="4" />
                <ENTRY entrytime="00:00:57.84" eventid="1277" heatid="40309" lane="8">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:00:58.29" />
                </ENTRY>
                <ENTRY entrytime="00:04:48.68" eventid="1073" heatid="40001" lane="5">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-14" qualificationtime="00:04:48.68" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Kim Sophie" lastname="Franke" birthdate="2013-01-01" gender="F" nation="GER" license="443664" athleteid="39670">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.92" eventid="1367" heatid="40445" lane="1">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:36.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.69" eventid="1227" heatid="40200" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:20.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.40" eventid="1123" heatid="40034" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:33.40" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Gruner" birthdate="2013-01-01" gender="F" nation="GER" license="443666" athleteid="39444">
              <ENTRIES>
                <ENTRY entrytime="00:03:00.98" eventid="1347" heatid="40405" lane="5" />
                <ENTRY entrytime="00:01:20.98" eventid="1267" heatid="40263" lane="7">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:32.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.98" eventid="1327" heatid="40379" lane="2">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:47.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.98" eventid="1123" heatid="40027" lane="3">
                  <MEETINFO name="Stadtmeisterschaft Dresden" city="Dresden" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:42.22" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.98" eventid="1227" heatid="40192" lane="5">
                  <MEETINFO name="Stadtmeisterschaft Dresden" city="Dresden" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:01:52.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.98" eventid="1207" heatid="40159" lane="5">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:48.20" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Zesewitz" birthdate="2010-01-01" gender="M" nation="GER" license="412733" athleteid="39701">
              <ENTRIES>
                <ENTRY entrytime="00:02:25.22" eventid="1173" heatid="40139" lane="4" />
                <ENTRY entrytime="00:02:19.66" eventid="1317" heatid="40376" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:16.80" />
                </ENTRY>
                <ENTRY entrytime="00:04:16.83" eventid="1257" heatid="40259" lane="5">
                  <MEETINFO name="136. Deutsche Meisterschaften im Schwimmen" city="Berlin" course="LCM" approved="GER" date="2025-05-01" qualificationtime="00:04:16.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.04" eventid="1357" heatid="40437" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:00.20" />
                </ENTRY>
                <ENTRY entrytime="00:04:45.97" eventid="1073" heatid="40002" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:04:44.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Max" lastname="Kolkowski" birthdate="2015-01-01" gender="M" nation="GER" license="463197" athleteid="39897">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.71" eventid="1217" heatid="40177" lane="1">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:44.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.45" eventid="1377" heatid="40462" lane="2">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:39.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.85" eventid="1297" heatid="40333" lane="2">
                  <MEETINFO name="Giraffenpokal" city="Chemnitz" course="LCM" approved="GER" date="2025-11-08" qualificationtime="00:00:37.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.61" eventid="1237" heatid="40218" lane="1">
                  <MEETINFO name="Giraffenpokal" city="Chemnitz" course="LCM" approved="GER" date="2025-11-08" qualificationtime="00:01:27.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.57" eventid="1337" heatid="40393" lane="7">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:37.57" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.64" eventid="1357" heatid="40423" lane="3">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:02:49.64" />
                </ENTRY>
                <ENTRY entrytime="00:03:34.86" eventid="1153" heatid="40102" lane="3">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:03:34.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Arian" lastname="Wüstenhagen" birthdate="2006-01-01" gender="M" nation="GER" license="349848" athleteid="39283">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.82" eventid="1337" heatid="40403" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:00.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.75" eventid="1397" heatid="40497" lane="7">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:55.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.44" eventid="1217" heatid="40190" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.25" eventid="1377" heatid="40473" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:26.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Elias" lastname="Conseur" birthdate="2015-01-01" gender="M" nation="GER" license="463192" athleteid="39805">
              <ENTRIES>
                <ENTRY entrytime="00:01:26.63" eventid="1237" heatid="40218" lane="5">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:26.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.84" eventid="1277" heatid="40291" lane="3">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:16.84" />
                </ENTRY>
                <ENTRY entrytime="00:03:09.78" eventid="1317" heatid="40364" lane="1">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:03:09.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.86" eventid="1217" heatid="40174" lane="1">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:49.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.65" eventid="1133" heatid="40063" lane="3">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:33.06" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.06" eventid="1173" heatid="40130" lane="3">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:03:05.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.68" eventid="1397" heatid="40487" lane="7">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:27.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nienke" lastname="Rudolph" birthdate="2014-01-01" gender="F" nation="GER" license="448172" athleteid="39553">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.76" eventid="1367" heatid="40447" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:37.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.72" eventid="1327" heatid="40386" lane="2">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:23.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.74" eventid="1207" heatid="40162" lane="1">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:41.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.01" eventid="1307" heatid="40356" lane="1">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:47.83" />
                </ENTRY>
                <ENTRY entrytime="00:03:16.46" eventid="1143" heatid="40093" lane="3">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:03:16.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.74" eventid="1123" heatid="40030" lane="3">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:33.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.39" eventid="1227" heatid="40200" lane="5">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:17.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Charlotte" lastname="Matthes" birthdate="2015-01-01" gender="F" nation="GER" license="463217" athleteid="39984">
              <ENTRIES>
                <ENTRY entrytime="00:12:00.00" eventid="1083" heatid="40004" lane="8" />
                <ENTRY entrytime="00:00:34.73" eventid="1123" heatid="40030" lane="5">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:33.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.23" eventid="1227" heatid="40197" lane="3">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:25.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.76" eventid="1267" heatid="40265" lane="3">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:01:17.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.41" eventid="1347" heatid="40407" lane="2">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:02:49.41" />
                </ENTRY>
                <ENTRY entrytime="00:03:04.15" eventid="1163" heatid="40115" lane="6">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:03:04.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.83" eventid="1367" heatid="40445" lane="2">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:37.82" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sirko" lastname="Sperling" birthdate="2014-01-01" gender="M" nation="GER" license="452436" athleteid="39780">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.39" eventid="1237" heatid="40223" lane="8">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:19.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.77" eventid="1217" heatid="40178" lane="7">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:39.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.04" eventid="1357" heatid="40424" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:45.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.77" eventid="1173" heatid="40131" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:59.77" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.33" eventid="1133" heatid="40068" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:31.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.42" eventid="1317" heatid="40367" lane="6">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:02:51.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.15" eventid="1337" heatid="40395" lane="3">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:30.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.00" eventid="1185" heatid="40146" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="39317" number="1" />
                    <RELAYPOSITION athleteid="39283" number="2" />
                    <RELAYPOSITION athleteid="39713" number="3" />
                    <RELAYPOSITION athleteid="39629" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" date="2025-10-26" qualificationtime="00:01:46.84" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.00" eventid="1185" heatid="40146" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" date="2025-10-26" qualificationtime="00:01:46.84" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:01:57.50" eventid="1183" heatid="40144" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" date="2025-10-26" qualificationtime="00:01:56.73" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <ENTRIES>
                <ENTRY entrytime="00:02:15.00" eventid="1183" heatid="40144" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" date="2025-10-26" qualificationtime="00:01:56.73" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5139" nation="GER" region="04" clubid="38790" name="SSV Senftenberg e.V.">
          <ATHLETES>
            <ATHLETE firstname="Martin" lastname="Schultz" birthdate="2009-01-01" gender="M" nation="GER" license="408377" athleteid="38834">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.52" eventid="1133" heatid="40077" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:28.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.95" eventid="1173" heatid="40138" lane="1">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:02:36.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.87" eventid="1217" heatid="40183" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:35.71" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.10" eventid="1237" heatid="40227" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:10.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.07" eventid="1277" heatid="40301" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:02.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.85" eventid="1297" heatid="40337" lane="3">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:32.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.22" eventid="1377" heatid="40470" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:32.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Edwin" lastname="Krosta" birthdate="2014-01-01" gender="M" nation="GER" license="490054" athleteid="38816">
              <ENTRIES>
                <ENTRY entrytime="00:01:29.99" eventid="1277" heatid="40287" lane="2">
                  <MEETINFO name="6. Frühjahrswettkampf" city="Dresden" course="SCM" approved="GER" date="2025-03-23" qualificationtime="00:01:38.29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="1297" heatid="40331" lane="7">
                  <MEETINFO name="Talentewettkampf" city="Cottbus" course="SCM" approved="GER" date="2025-06-22" qualificationtime="00:01:07.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:48.99" eventid="1377" heatid="40460" lane="6">
                  <MEETINFO name="6. Frühjahrswettkampf" city="Dresden" course="SCM" approved="GER" date="2025-03-23" qualificationtime="00:00:54.45" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Rebecca" lastname="Hoffmann" birthdate="2015-01-01" gender="F" nation="GER" license="448398" athleteid="38800">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.62" eventid="1123" heatid="40029" lane="2">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:35.62" />
                </ENTRY>
                <ENTRY entrytime="00:03:14.42" eventid="1163" heatid="40113" lane="5">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:03:14.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.04" eventid="1207" heatid="40157" lane="3">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:56.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.43" eventid="1227" heatid="40192" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:32.95" />
                </ENTRY>
                <ENTRY entrytime="00:07:21.40" eventid="1247" heatid="40233" lane="3">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:07:21.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.78" eventid="1267" heatid="40264" lane="1">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:17.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.26" eventid="1287" heatid="40313" lane="2">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:39.26" />
                </ENTRY>
                <ENTRY entrytime="00:03:31.99" eventid="1307" heatid="40348" lane="2">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:03:21.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.84" eventid="1347" heatid="40406" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:57.16" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.11" eventid="1367" heatid="40441" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:42.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.27" eventid="1387" heatid="40475" lane="3">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:28.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Maurer" birthdate="2009-01-01" gender="F" nation="GER" license="453444" athleteid="38824">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.41" eventid="1123" heatid="40037" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:31.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.31" eventid="1267" heatid="40272" lane="3">
                  <MEETINFO name="Double-Pool-Meeting (25m Bahn)" city="Riesa" course="SCM" approved="GER" date="2025-02-08" qualificationtime="00:01:10.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Charly" lastname="Krosta" birthdate="2014-01-01" gender="M" nation="GER" license="490055" athleteid="38812">
              <ENTRIES>
                <ENTRY entrytime="00:01:28.99" eventid="1277" heatid="40287" lane="6">
                  <MEETINFO name="6. Frühjahrswettkampf" city="Dresden" course="SCM" approved="GER" date="2025-03-23" qualificationtime="00:01:32.89" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="1297" heatid="40331" lane="6">
                  <MEETINFO name="36. Lagen – Srintpokal des SSV Senftenberg e.V." city="Senftenberg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:50.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:48.99" eventid="1377" heatid="40460" lane="3">
                  <MEETINFO name="31. Delphinpokal" city="Ludwigsfelde" course="SCM" approved="GER" date="2025-01-18" qualificationtime="00:00:48.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Oliver" lastname="Hoffmann" birthdate="2011-01-01" gender="M" nation="GER" license="408376" athleteid="38791">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.01" eventid="1133" heatid="40076" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:28.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.84" eventid="1237" heatid="40222" lane="5">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:01:19.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.82" eventid="1277" heatid="40299" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:05.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.82" eventid="1297" heatid="40338" lane="8">
                  <MEETINFO name="31. Delphinpokal" city="Ludwigsfelde" course="SCM" approved="GER" date="2025-01-18" qualificationtime="00:00:31.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.49" eventid="1317" heatid="40368" lane="3">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:02:48.49" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.65" eventid="1357" heatid="40425" lane="3">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:02:36.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.40" eventid="1377" heatid="40468" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:34.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.04" eventid="1397" heatid="40490" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:15.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Timo" lastname="Schorten" birthdate="2008-01-01" gender="M" nation="GER" license="446904" athleteid="38827">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.57" eventid="1133" heatid="40081" lane="8">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:00:27.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.15" eventid="1277" heatid="40303" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:02.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.14" eventid="1297" heatid="40343" lane="1">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:28.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.24" eventid="1357" heatid="40431" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:20.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.49" eventid="1377" heatid="40469" lane="5">
                  <MEETINFO name="36. Lagen – Srintpokal des SSV Senftenberg e.V." city="Senftenberg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:31.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.92" eventid="1397" heatid="40492" lane="4">
                  <MEETINFO name="Offene Thüringer Meisterschaften" city="Erfurt" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:07.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Manuel" lastname="Lehning" birthdate="2013-01-01" gender="M" nation="GER" license="490056" athleteid="38820">
              <ENTRIES>
                <ENTRY entrytime="00:01:25.99" eventid="1277" heatid="40288" lane="1">
                  <MEETINFO name="36. Lagen – Srintpokal des SSV Senftenberg e.V." city="Senftenberg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:38.21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="1297" heatid="40331" lane="2" />
                <ENTRY entrytime="00:00:44.99" eventid="1377" heatid="40461" lane="1">
                  <MEETINFO name="36. Lagen – Srintpokal des SSV Senftenberg e.V." city="Senftenberg" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:49.84" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Luise" lastname="Thieß" birthdate="2009-01-01" gender="F" nation="GER" license="379286" athleteid="38842">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.55" eventid="1287" heatid="40319" lane="8">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:00:35.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.03" eventid="1367" heatid="40451" lane="1">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:00:37.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Hendrik" gender="M" lastname="Just" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="6506" nation="GER" region="12" clubid="38483" name="Schwimmsportverein Kirschau e.V.">
          <ATHLETES>
            <ATHLETE firstname="Fabio" lastname="Gerber" birthdate="2007-01-01" gender="M" nation="GER" license="397578" athleteid="38490">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.45" eventid="1133" heatid="40081" lane="1">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:26.02" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.85" eventid="1153" heatid="40107" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:58.85" />
                </ENTRY>
                <ENTRY entrytime="00:04:40.00" eventid="1257" heatid="40257" lane="3" />
                <ENTRY entrytime="00:01:00.02" eventid="1277" heatid="40306" lane="8">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:01:00.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.47" eventid="1297" heatid="40341" lane="8">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:00:29.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.00" eventid="1317" heatid="40373" lane="8" />
                <ENTRY entrytime="00:01:17.71" eventid="1337" heatid="40400" lane="6">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:01:13.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.49" eventid="1357" heatid="40433" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:14.49" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Jannasch" birthdate="2012-01-01" gender="M" nation="GER" license="484093" athleteid="38507">
              <ENTRIES>
                <ENTRY entrytime="00:10:45.00" eventid="1093" heatid="40014" lane="2" />
                <ENTRY entrytime="00:00:36.80" eventid="1133" heatid="40061" lane="7">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:00:36.80" />
                </ENTRY>
                <ENTRY entrytime="00:03:25.00" eventid="1153" heatid="40103" lane="6" />
                <ENTRY entrytime="00:01:27.00" eventid="1237" heatid="40218" lane="2" />
                <ENTRY entrytime="00:05:10.00" eventid="1257" heatid="40253" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Charly" lastname="Reinsch" birthdate="2015-01-01" gender="M" nation="GER" license="499558" athleteid="38526">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.41" eventid="1133" heatid="40059" lane="3">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:00:41.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.53" eventid="1217" heatid="40174" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:00:54.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.87" eventid="1377" heatid="40460" lane="2">
                  <MEETINFO name="EnjoyQuality Bonbon Pokal" city="Zittau" course="SCM" approved="GER" date="2025-03-15" qualificationtime="00:00:50.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nikolas" lastname="Kühnel" birthdate="2010-01-01" gender="M" nation="GER" license="469955" athleteid="38517">
              <ENTRIES>
                <ENTRY entrytime="00:02:59.00" eventid="1153" heatid="40106" lane="4" />
                <ENTRY entrytime="00:00:37.08" eventid="1217" heatid="40183" lane="8">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:36.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.24" eventid="1297" heatid="40335" lane="1">
                  <MEETINFO name="Frühjahrsschwimmfest" city="Görlitz" course="SCM" approved="GER" date="2025-03-29" qualificationtime="00:00:34.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.87" eventid="1337" heatid="40398" lane="8">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:01:21.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alina" lastname="Hnatchenko" birthdate="2011-01-01" gender="F" nation="UKR" license="463688" athleteid="38499">
              <ENTRIES>
                <ENTRY entrytime="00:11:20.00" eventid="1083" heatid="40006" lane="1" />
                <ENTRY entrytime="00:00:34.26" eventid="1123" heatid="40031" lane="4">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:00:33.66" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.61" eventid="1163" heatid="40114" lane="2">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:03:07.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.43" eventid="1227" heatid="40196" lane="2">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:01:24.89" />
                </ENTRY>
                <ENTRY entrytime="00:05:19.00" eventid="1247" heatid="40239" lane="5" />
                <ENTRY entrytime="00:01:15.69" eventid="1267" heatid="40266" lane="5">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:01:15.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.08" eventid="1367" heatid="40442" lane="4">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:38.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Bennet" lastname="Brock" birthdate="2010-01-01" gender="M" nation="GER" license="430118" athleteid="38484">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.29" eventid="1133" heatid="40078" lane="3">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:00:27.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.00" eventid="1237" heatid="40223" lane="2" />
                <ENTRY entrytime="00:01:03.37" eventid="1277" heatid="40301" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:03.37" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.89" eventid="1297" heatid="40339" lane="2">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:00:31.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.26" eventid="1377" heatid="40468" lane="2">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:00:33.70" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Schmidt" birthdate="2009-01-01" gender="M" nation="GER" license="510041" athleteid="38540">
              <ENTRIES>
                <ENTRY entrytime="00:04:39.00" eventid="1257" heatid="40258" lane="1" />
                <ENTRY entrytime="00:01:02.00" eventid="1277" heatid="40303" lane="6">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:01:09.70" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lotta" lastname="Jannasch" birthdate="2014-01-01" gender="F" nation="GER" license="469951" athleteid="38513">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.66" eventid="1123" heatid="40026" lane="7">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:00:40.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.18" eventid="1207" heatid="40157" lane="5">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:00:55.18" />
                </ENTRY>
                <ENTRY entrytime="00:06:00.00" eventid="1247" heatid="40235" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Frederic" lastname="Nehrettig" birthdate="2009-01-01" gender="M" nation="GER" license="440166" athleteid="38522">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.89" eventid="1133" heatid="40073" lane="7">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:29.78" />
                </ENTRY>
                <ENTRY entrytime="00:04:40.00" eventid="1257" heatid="40257" lane="4" />
                <ENTRY entrytime="00:01:08.49" eventid="1277" heatid="40297" lane="7">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:01:07.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leonie" lastname="Schierz" birthdate="2012-01-01" gender="F" nation="GER" license="463589" athleteid="38530">
              <ENTRIES>
                <ENTRY entrytime="00:11:20.00" eventid="1083" heatid="40006" lane="7" />
                <ENTRY entrytime="00:00:35.74" eventid="1123" heatid="40028" lane="4">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:00:34.20" />
                </ENTRY>
                <ENTRY entrytime="00:03:25.00" eventid="1143" heatid="40092" lane="8" />
                <ENTRY entrytime="00:00:43.80" eventid="1207" heatid="40160" lane="3">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:43.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.99" eventid="1227" heatid="40196" lane="8">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:01:27.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.65" eventid="1267" heatid="40264" lane="7">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:01:14.27" />
                </ENTRY>
                <ENTRY entrytime="00:03:09.00" eventid="1307" heatid="40349" lane="5" />
                <ENTRY entrytime="00:01:38.97" eventid="1327" heatid="40379" lane="4">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:01:33.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.88" eventid="1367" heatid="40443" lane="7">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:37.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.00" eventid="1185" heatid="40146" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="38490" number="1" />
                    <RELAYPOSITION athleteid="38522" number="2" />
                    <RELAYPOSITION athleteid="38540" number="3" />
                    <RELAYPOSITION athleteid="38507" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="3410" nation="GER" region="12" clubid="38259" name="USV TU Dresden e.V.">
          <ATHLETES>
            <ATHLETE firstname="Jonas" lastname="Kuhtz" birthdate="2010-01-01" gender="M" nation="GER" license="441838" athleteid="38307">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.20" eventid="1133" heatid="40079" lane="8">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:27.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.63" eventid="1297" heatid="40338" lane="7">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:31.77" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.75" eventid="1377" heatid="40472" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:29.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.18" eventid="1173" heatid="40136" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:32.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.26" eventid="1217" heatid="40183" lane="5">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:35.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hugo" lastname="Schütze" birthdate="2011-01-01" gender="M" nation="GER" license="426686" athleteid="38376">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.26" eventid="1133" heatid="40078" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:27.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.22" eventid="1217" heatid="40184" lane="8">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:36.22" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.97" eventid="1277" heatid="40303" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:01.49" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.83" eventid="1337" heatid="40398" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:16.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.84" eventid="1357" heatid="40430" lane="3">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:02:19.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Kirill" lastname="Kurlykov" birthdate="2012-01-01" gender="M" nation="GER" license="437629" athleteid="38313">
              <ENTRIES>
                <ENTRY entrytime="00:02:22.78" eventid="1357" heatid="40430" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:21.45" />
                </ENTRY>
                <ENTRY entrytime="00:05:48.00" eventid="1073" heatid="39999" lane="5">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-26" qualificationtime="00:05:48.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.51" eventid="1317" heatid="40371" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:37.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.51" eventid="1277" heatid="40299" lane="7">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:01:05.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.86" eventid="1133" heatid="40073" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:29.23" />
                </ENTRY>
                <ENTRY entrytime="00:05:07.04" eventid="1257" heatid="40253" lane="5">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:05:07.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.99" eventid="1237" heatid="40226" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:01:13.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Max" lastname="Schwarzer" birthdate="2011-01-01" gender="M" nation="GER" license="437639" athleteid="38382">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.38" eventid="1133" heatid="40070" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:31.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.84" eventid="1237" heatid="40221" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:16.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.84" eventid="1277" heatid="40294" lane="5">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:08.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.02" eventid="1297" heatid="40335" lane="3">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:34.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.50" eventid="1377" heatid="40465" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:35.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jonas" lastname="Langner" birthdate="2009-01-01" gender="M" nation="GER" license="395538" athleteid="38321">
              <ENTRIES>
                <ENTRY entrytime="00:02:26.43" eventid="1317" heatid="40373" lane="3">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:02:26.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.33" eventid="1133" heatid="40081" lane="3">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:26.69" />
                </ENTRY>
                <ENTRY entrytime="00:09:09.83" eventid="1093" heatid="40018" lane="4">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:09:09.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.90" eventid="1357" heatid="40435" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:04.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Tilman" lastname="Sachs" birthdate="2001-01-01" gender="M" nation="GER" license="249621" athleteid="38360">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.86" eventid="1133" heatid="40088" lane="2">
                  <MEETINFO name="Double-Pool-Meeting (25m Bahn)" city="Riesa" course="SCM" approved="GER" date="2025-02-08" qualificationtime="00:00:24.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.02" eventid="1217" heatid="40189" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:29.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.07" eventid="1277" heatid="40310" lane="4">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:54.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.31" eventid="1337" heatid="40403" lane="8">
                  <MEETINFO name="28. DMSM Bundesentscheid" city="Nürnberg" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:03.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maik" lastname="Punke" birthdate="1997-01-01" gender="M" nation="GER" license="392584" athleteid="38348">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.37" eventid="1133" heatid="40085" lane="1">
                  <MEETINFO name="Starker August" city="Dresden" course="LCM" approved="GER" date="2025-02-01" qualificationtime="00:00:26.37" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.62" eventid="1217" heatid="40188" lane="5">
                  <MEETINFO name="Deutsche Hochschulmeisterschaft Schwimmen" city="Düsseldorf" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:31.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Dittel" birthdate="2012-01-01" gender="F" nation="GER" license="437623" athleteid="38260">
              <ENTRIES>
                <ENTRY entrytime="00:10:23.91" eventid="1083" heatid="40009" lane="4">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:10:23.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.75" eventid="1163" heatid="40127" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:24.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.16" eventid="1347" heatid="40418" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:13.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.45" eventid="1227" heatid="40212" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:07.31" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.61" eventid="1267" heatid="40284" lane="8">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:01:02.61" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.16" eventid="1367" heatid="40458" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:31.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.81" eventid="1307" heatid="40358" lane="6">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:39.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sascha" lastname="Grams" birthdate="2015-01-01" gender="M" nation="GER" license="471326" athleteid="38290">
              <ENTRIES>
                <ENTRY entrytime="00:06:13.07" eventid="1257" heatid="40246" lane="3">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:06:13.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.66" eventid="1217" heatid="40176" lane="2">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:44.03" />
                </ENTRY>
                <ENTRY entrytime="00:04:17.62" eventid="1153" heatid="40101" lane="3">
                  <MEETINFO name="Stadtmeisterschaft Dresden" city="Dresden" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:04:17.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:39.72" eventid="1337" heatid="40393" lane="8">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:01:39.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.77" eventid="1277" heatid="40292" lane="5">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:14.46" />
                </ENTRY>
                <ENTRY entrytime="00:03:15.26" eventid="1317" heatid="40363" lane="7">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:03:04.27" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leonard" lastname="Tkachenko" birthdate="2010-01-01" gender="M" nation="GER" license="410656" athleteid="38395">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.82" eventid="1133" heatid="40071" lane="2">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:29.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.74" eventid="1217" heatid="40182" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:37.74" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Eisert" birthdate="2012-01-01" gender="F" nation="GER" license="437624" athleteid="38274">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.20" eventid="1123" heatid="40049" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:29.98" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.55" eventid="1227" heatid="40204" lane="3">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:14.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.20" eventid="1267" heatid="40278" lane="5">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:05.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.43" eventid="1347" heatid="40414" lane="3">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:02:28.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.95" eventid="1367" heatid="40451" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:34.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anton" lastname="Sukhanov" birthdate="2006-01-01" gender="M" nation="GER" license="336098" athleteid="38390">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.00" eventid="1133" heatid="40083" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:27.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.70" eventid="1217" heatid="40187" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:32.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.63" eventid="1297" heatid="40342" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:28.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.77" eventid="1337" heatid="40400" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:11.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Franziska" lastname="Grammlich" birthdate="2005-01-01" gender="F" nation="GER" license="349778" athleteid="38280">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.92" eventid="1227" heatid="40213" lane="2">
                  <MEETINFO name="DMSM Berlin" city="Berlin" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:06.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.42" eventid="1367" heatid="40459" lane="7">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-30" qualificationtime="00:00:32.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.63" eventid="1267" heatid="40285" lane="4">
                  <MEETINFO name="DMSM Berlin" city="Berlin" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:00.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lukas" lastname="Langner" birthdate="2011-01-01" gender="M" nation="GER" license="426678" athleteid="38326">
              <ENTRIES>
                <ENTRY entrytime="00:02:28.27" eventid="1317" heatid="40373" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:28.27" />
                </ENTRY>
                <ENTRY entrytime="00:09:25.03" eventid="1093" heatid="40018" lane="6">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:09:25.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.57" eventid="1133" heatid="40077" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:28.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.95" eventid="1277" heatid="40303" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:00.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.20" eventid="1377" heatid="40472" lane="8">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:31.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.93" eventid="1237" heatid="40230" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:05.49" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.53" eventid="1173" heatid="40139" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:18.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Katharina" lastname="Grammlich" birthdate="2008-01-01" gender="F" nation="GER" license="380800" athleteid="38284">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.38" eventid="1367" heatid="40459" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:30.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.53" eventid="1163" heatid="40127" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:24.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.19" eventid="1307" heatid="40358" lane="1" />
                <ENTRY entrytime="00:00:29.35" eventid="1123" heatid="40053" lane="6" />
                <ENTRY entrytime="00:01:08.43" eventid="1227" heatid="40213" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:05.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ella" lastname="Schumann" birthdate="2011-01-01" gender="F" nation="GER" license="426684" athleteid="38365">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.30" eventid="1123" heatid="40038" lane="1">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:00:32.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.28" eventid="1227" heatid="40201" lane="8">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:19.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.71" eventid="1267" heatid="40268" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:13.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.64" eventid="1287" heatid="40315" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:36.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.44" eventid="1367" heatid="40446" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:36.67" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Keusch" birthdate="1995-01-01" gender="F" nation="GER" license="172579" athleteid="38303">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.41" eventid="1123" heatid="40048" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:30.41" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.00" eventid="1163" heatid="40119" lane="5">
                  <MEETINFO name="39. Internationale DM Masters Lange Strecke" city="Wolfsburg" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:02:49.20" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.00" eventid="1247" heatid="40241" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:05:14.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Theresa" lastname="Einbock" birthdate="2012-01-01" gender="F" nation="GER" license="445207" athleteid="38268">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.20" eventid="1123" heatid="40038" lane="3">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:00:32.20" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.99" eventid="1207" heatid="40170" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:37.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.66" eventid="1267" heatid="40269" lane="5">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:11.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.85" eventid="1287" heatid="40324" lane="8">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:00:32.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.07" eventid="1327" heatid="40388" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:23.07" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Moritz" lastname="Jacob" birthdate="2010-01-01" gender="M" nation="GER" license="410639" athleteid="38297">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.43" eventid="1133" heatid="40075" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:28.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.69" eventid="1277" heatid="40300" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:01.16" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.06" eventid="1297" heatid="40339" lane="8">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:00:32.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.89" eventid="1357" heatid="40429" lane="7">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:02:22.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.19" eventid="1377" heatid="40468" lane="3">
                  <MEETINFO name="14. Sängerpokal" city="Finsterwalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:00:33.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lea-Sophie" lastname="Maihold" birthdate="2011-01-01" gender="F" nation="GER" license="437630" athleteid="38334">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.45" eventid="1123" heatid="40044" lane="1">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:30.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.92" eventid="1207" heatid="40163" lane="2">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:41.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.60" eventid="1267" heatid="40276" lane="2">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:07.61" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.94" eventid="1307" heatid="40354" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:02:53.94" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.51" eventid="1347" heatid="40412" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:02:34.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nico" lastname="Stechemesser" birthdate="1975-01-01" gender="M" nation="GER" license="128152" athleteid="38388">
              <ENTRIES>
                <ENTRY entrytime="00:21:21.21" eventid="1113" heatid="40023" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alexander" lastname="Paulin" birthdate="2004-01-01" gender="M" nation="GER" license="315754" athleteid="38343">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.43" eventid="1133" heatid="40084" lane="4">
                  <MEETINFO name="TuR´s Hexentanz" city="Dresden" course="SCM" approved="GER" date="2025-04-26" qualificationtime="00:00:26.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.78" eventid="1277" heatid="40304" lane="5">
                  <MEETINFO name="TuR´s Hexentanz" city="Dresden" course="SCM" approved="GER" date="2025-04-26" qualificationtime="00:01:00.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.50" eventid="1297" heatid="40344" lane="1">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-30" qualificationtime="00:00:28.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.30" eventid="1397" heatid="40492" lane="7">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:01:07.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lukas" lastname="Ranft" birthdate="2011-01-01" gender="M" nation="GER" license="426681" athleteid="38351">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.53" eventid="1133" heatid="40077" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:28.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.47" eventid="1217" heatid="40180" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:36.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Mehrholz" birthdate="1974-01-01" gender="M" nation="GER" license="444423" athleteid="38340">
              <ENTRIES>
                <ENTRY entrytime="00:18:30.00" eventid="1113" status="WDR" heatid="40025" lane="6" />
                <ENTRY entrytime="00:00:27.00" eventid="1133" status="WDR" heatid="40083" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:27.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Margot" lastname="Schumann" birthdate="2012-01-01" gender="F" nation="GER" license="437638" athleteid="38371">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.13" eventid="1123" heatid="40029" lane="5">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:34.96" />
                </ENTRY>
                <ENTRY entrytime="00:03:26.93" eventid="1143" heatid="40091" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:03:10.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.73" eventid="1207" heatid="40165" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:39.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.06" eventid="1327" heatid="40382" lane="4">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:27.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Henriette" lastname="Rex" birthdate="2011-01-01" gender="F" nation="GER" license="426682" athleteid="38354">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.72" eventid="1123" heatid="40042" lane="3">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:00:31.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.25" eventid="1227" heatid="40198" lane="6">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:18.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.24" eventid="1267" heatid="40271" lane="7">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:09.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.37" eventid="1347" heatid="40409" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:39.37" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.56" eventid="1367" heatid="40446" lane="1">
                  <MEETINFO name="14. Sängerpokal" city="Finsterwalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:00:37.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3603" nation="GER" region="13" clubid="38622" name="SSV 70 Halle-Neustadt">
          <ATHLETES>
            <ATHLETE firstname="Niklas" lastname="Rüssel" birthdate="2014-01-01" gender="M" nation="GER" license="464816" athleteid="38728">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.60" eventid="1133" heatid="40065" lane="2">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:33.60" />
                </ENTRY>
                <ENTRY entrytime="00:03:33.15" eventid="1153" heatid="40102" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:33.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.33" eventid="1217" heatid="40178" lane="8">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:43.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.94" eventid="1237" heatid="40218" lane="6">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:26.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.03" eventid="1277" heatid="40293" lane="1">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:01:15.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.32" eventid="1337" heatid="40394" lane="1">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:34.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leah Sophie" lastname="Bauer" birthdate="2010-01-01" gender="F" nation="GER" license="406166" athleteid="38623">
              <ENTRIES>
                <ENTRY entrytime="00:02:36.82" eventid="1163" heatid="40125" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:02:30.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.12" eventid="1227" heatid="40212" lane="6">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:01:08.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.04" eventid="1307" heatid="40358" lane="8" />
                <ENTRY entrytime="00:00:32.45" eventid="1367" heatid="40458" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:31.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Klausnitz" birthdate="2014-01-01" gender="M" nation="GER" license="452347" athleteid="38686">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.71" eventid="1133" heatid="40067" lane="6">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:32.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.41" eventid="1173" heatid="40132" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:56.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.38" eventid="1237" heatid="40224" lane="1">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:17.38" />
                </ENTRY>
                <ENTRY entrytime="00:05:31.74" eventid="1257" heatid="40249" lane="2">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:05:31.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.50" eventid="1277" heatid="40296" lane="3">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:09.50" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.16" eventid="1317" heatid="40367" lane="1">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:53.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Sachadae" birthdate="2011-01-01" gender="M" nation="GER" license="427208" athleteid="38735">
              <ENTRIES>
                <ENTRY entrytime="00:18:46.87" eventid="1113" heatid="40025" lane="7" />
                <ENTRY entrytime="00:02:18.83" eventid="1197" heatid="40156" lane="8">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:02:15.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.90" eventid="1237" heatid="40230" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:01.90" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.07" eventid="1277" heatid="40309" lane="3">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:54.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.75" eventid="1397" heatid="40496" lane="6">
                  <MEETINFO name="30. Norddeutscher Jugendländervergleich" city="Lübeck" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:01:00.52" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Julius" lastname="Luci" birthdate="2008-01-01" gender="M" nation="GER" license="391868" athleteid="38697">
              <ENTRIES>
                <ENTRY entrytime="00:02:39.89" eventid="1153" heatid="40110" lane="2">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:02:39.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.77" eventid="1217" heatid="40187" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:31.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.88" eventid="1317" heatid="40376" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:19.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.53" eventid="1397" heatid="40494" lane="2">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:02.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Wolff" birthdate="2009-01-01" gender="M" nation="GER" license="409316" athleteid="38764">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.13" eventid="1133" heatid="40085" lane="3">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:25.79" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.46" eventid="1237" heatid="40229" lane="6">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:06.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.83" eventid="1277" heatid="40307" lane="5">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:57.04" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.16" eventid="1357" heatid="40435" lane="5">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:02:06.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emma Leni" lastname="Schulz" birthdate="2014-01-01" gender="F" nation="GER" license="450929" athleteid="38746">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.23" eventid="1123" heatid="40038" lane="6">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:32.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.06" eventid="1163" heatid="40119" lane="1">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:51.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.30" eventid="1227" heatid="40205" lane="5">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:17.30" />
                </ENTRY>
                <ENTRY entrytime="00:05:24.85" eventid="1247" heatid="40238" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:05:24.85" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.94" eventid="1307" heatid="40356" lane="6">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:48.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.51" eventid="1327" heatid="40382" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lotta" lastname="Hanning" birthdate="2009-01-01" gender="F" nation="GER" license="396628" athleteid="38663">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.97" eventid="1123" heatid="40046" lane="2">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:30.96" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.17" eventid="1163" heatid="40121" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:45.17" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.08" eventid="1227" heatid="40207" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:14.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.21" eventid="1267" heatid="40275" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:08.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.53" eventid="1367" heatid="40452" lane="7">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:34.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alexandra" lastname="Rennefahrt" birthdate="2008-01-01" gender="F" nation="GER" license="391869" athleteid="38716">
              <ENTRIES>
                <ENTRY entrytime="00:02:38.41" eventid="1163" heatid="40124" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:39.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.87" eventid="1207" heatid="40172" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:35.77" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.22" eventid="1327" heatid="40390" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:16.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.00" eventid="1367" heatid="40455" lane="5">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:34.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jakob" lastname="Rüssel" birthdate="2014-01-01" gender="M" nation="GER" license="464815" athleteid="38721">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.16" eventid="1133" heatid="40062" lane="4">
                  <MEETINFO name="Kids-Cup Teil 1 des LSVSA der Leistungsstützpunkte" city="Bitterfeld-Wolfen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:35.16" />
                </ENTRY>
                <ENTRY entrytime="00:03:14.59" eventid="1173" heatid="40129" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:14.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.76" eventid="1217" heatid="40175" lane="7">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:47.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.45" eventid="1237" heatid="40216" lane="6">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:31.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.43" eventid="1277" heatid="40290" lane="7">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:01:19.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.99" eventid="1297" heatid="40332" lane="3">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:39.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Carl" lastname="Ertle" birthdate="2011-01-01" gender="M" nation="GER" license="436530" athleteid="38645">
              <ENTRIES>
                <ENTRY entrytime="00:02:54.78" eventid="1153" heatid="40108" lane="8">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:54.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.21" eventid="1237" heatid="40229" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:06.73" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.97" eventid="1317" heatid="40372" lane="2">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:34.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.65" eventid="1397" heatid="40492" lane="6">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:08.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Felsch" birthdate="2012-01-01" gender="F" nation="GER" license="436522" athleteid="38650">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.13" eventid="1207" heatid="40170" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:38.14" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.62" eventid="1227" heatid="40200" lane="3">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:01:22.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.31" eventid="1287" heatid="40322" lane="2">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:32.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.74" eventid="1367" heatid="40454" lane="1">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:00:34.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.65" eventid="1387" heatid="40481" lane="5">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:01:11.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Luzie" lastname="Petzold" birthdate="2013-01-01" gender="F" nation="GER" license="450925" athleteid="38709">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.62" eventid="1123" heatid="40036" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:32.62" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.29" eventid="1163" heatid="40115" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:03.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.23" eventid="1227" heatid="40206" lane="1">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:17.23" />
                </ENTRY>
                <ENTRY entrytime="00:05:46.59" eventid="1247" heatid="40236" lane="1">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:05:46.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.63" eventid="1267" heatid="40276" lane="7">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:08.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.61" eventid="1307" heatid="40352" lane="7">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:58.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Finn" lastname="Kochmann" birthdate="2006-01-01" gender="M" nation="GER" license="351810" athleteid="38693">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.89" eventid="1277" heatid="40311" lane="1" />
                <ENTRY entrytime="00:00:26.99" eventid="1297" heatid="40346" lane="2" />
                <ENTRY entrytime="00:00:28.65" eventid="1377" heatid="40473" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Elise" lastname="Zinnert" birthdate="2012-01-01" gender="F" nation="GER" license="436528" athleteid="38769">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.48" eventid="1123" heatid="40048" lane="2">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:30.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.46" eventid="1207" heatid="40169" lane="6">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:00:38.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.60" eventid="1267" heatid="40278" lane="1">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:04.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.50" eventid="1327" heatid="40387" lane="5">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:20.68" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.61" eventid="1347" heatid="40414" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:02:23.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nele" lastname="Behnert" birthdate="2011-01-01" gender="F" nation="GER" license="436526" athleteid="38628">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.40" eventid="1207" heatid="40164" lane="1">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:41.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.28" eventid="1227" heatid="40205" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:12.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.37" eventid="1327" heatid="40383" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:25.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.47" eventid="1367" heatid="40452" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:34.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Greta" lastname="Sosinski" birthdate="2011-01-01" gender="F" nation="GER" license="419503" athleteid="38753">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.01" eventid="1123" heatid="40055" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:28.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.41" eventid="1207" heatid="40167" lane="4" />
                <ENTRY entrytime="00:01:03.12" eventid="1267" heatid="40283" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:01.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.76" eventid="1307" heatid="40360" lane="8">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:02:34.76" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leni" lastname="Kehler" birthdate="2014-01-01" gender="F" nation="GER" license="450924" athleteid="38680">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.46" eventid="1123" heatid="40043" lane="4">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:31.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.37" eventid="1267" heatid="40278" lane="2">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:07.11" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.05" eventid="1307" heatid="40356" lane="8">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:02:46.77" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.58" eventid="1347" heatid="40415" lane="5">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:02:27.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.16" eventid="1387" heatid="40480" lane="7">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:15.40" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Evgenia" lastname="Bruch" birthdate="2010-01-01" gender="F" nation="GER" license="409314" athleteid="38639">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.08" eventid="1123" heatid="40054" lane="4">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:28.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.82" eventid="1227" heatid="40205" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:14.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.19" eventid="1267" heatid="40279" lane="2">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:04.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.98" eventid="1287" heatid="40323" lane="5">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:32.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.32" eventid="1367" heatid="40453" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:34.55" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Gutschlich" birthdate="2015-01-01" gender="F" nation="GER" license="464813" athleteid="38656">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.62" eventid="1123" heatid="40029" lane="7">
                  <MEETINFO name="Kids-Cup Teil 1 des LSVSA der Leistungsstützpunkte" city="Bitterfeld-Wolfen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:35.62" />
                </ENTRY>
                <ENTRY entrytime="00:03:32.59" eventid="1143" heatid="40091" lane="8">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:32.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.30" eventid="1207" heatid="40159" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:45.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.53" eventid="1227" heatid="40193" lane="8">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:01:35.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.44" eventid="1267" heatid="40264" lane="6">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:01:19.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.92" eventid="1327" heatid="40381" lane="1">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:34.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marisa Elin" lastname="Wilczek" birthdate="2009-01-01" gender="F" nation="GER" license="409308" athleteid="38758">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.54" eventid="1123" heatid="40052" lane="5">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:29.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.92" eventid="1227" heatid="40208" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:11.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.99" eventid="1267" heatid="40279" lane="4">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:04.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.69" eventid="1287" heatid="40324" lane="6">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:31.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.90" eventid="1367" heatid="40456" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:32.93" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Höllger" birthdate="2014-01-01" gender="F" nation="GER" license="450923" athleteid="38669">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.62" eventid="1143" heatid="40094" lane="6">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:03:09.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.35" eventid="1207" heatid="40164" lane="2">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:39.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.64" eventid="1287" heatid="40313" lane="8">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:00:39.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.15" eventid="1327" heatid="40384" lane="1">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:28.35" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jannik" lastname="Zorn" birthdate="2013-01-01" gender="M" nation="GER" license="450934" athleteid="38775">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.33" eventid="1133" heatid="40068" lane="2">
                  <MEETINFO name="Kids-Cup Teil 1 des LSVSA der Leistungsstützpunkte" city="Bitterfeld-Wolfen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:32.33" />
                </ENTRY>
                <ENTRY entrytime="00:03:11.78" eventid="1153" heatid="40105" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:03:11.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.91" eventid="1217" heatid="40179" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:41.91" />
                </ENTRY>
                <ENTRY entrytime="00:05:26.86" eventid="1257" heatid="40250" lane="6">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:05:26.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.65" eventid="1277" heatid="40297" lane="8">
                  <MEETINFO name="DMSJ" city="Burg" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:08.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.89" eventid="1337" heatid="40397" lane="6">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:22.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jan Henrik" lastname="Höllger" birthdate="2008-01-01" gender="M" nation="GER" license="391867" athleteid="38674">
              <ENTRIES>
                <ENTRY entrytime="00:18:07.44" eventid="1113" heatid="40025" lane="3" />
                <ENTRY entrytime="00:02:18.66" eventid="1197" heatid="40156" lane="1">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:02:16.53" />
                </ENTRY>
                <ENTRY entrytime="00:04:31.80" eventid="1257" heatid="40258" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:04:31.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.52" eventid="1297" heatid="40345" lane="7">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:27.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.95" eventid="1397" heatid="40496" lane="2">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:00.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fabian" lastname="Schalle" birthdate="2011-01-01" gender="M" nation="GER" license="436532" athleteid="38741">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.94" eventid="1133" heatid="40079" lane="5">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:27.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.11" eventid="1197" heatid="40153" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:45.11" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.57" eventid="1277" heatid="40302" lane="4">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:02.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.81" eventid="1397" heatid="40493" lane="3">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:01:06.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karl" lastname="Bönicke" birthdate="2013-01-01" gender="M" nation="GER" license="443919" athleteid="38633">
              <ENTRIES>
                <ENTRY entrytime="00:03:15.69" eventid="1153" heatid="40104" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:15.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.86" eventid="1173" heatid="40133" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:53.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.90" eventid="1237" heatid="40222" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:19.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:57.57" eventid="1317" heatid="40366" lane="7">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:02:57.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.95" eventid="1377" heatid="40464" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:36.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Luca" lastname="Mitrenga" birthdate="2008-01-01" gender="M" nation="GER" license="380826" athleteid="38702">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.70" eventid="1133" heatid="40087" lane="8">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:24.72" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.74" eventid="1173" heatid="40141" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:23.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.14" eventid="1237" heatid="40232" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:58.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.69" eventid="1297" heatid="40346" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:25.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.46" eventid="1317" heatid="40374" lane="2">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:02:23.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.00" eventid="1377" heatid="40474" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:27.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5274" nation="GER" region="14" clubid="34866" name="TSV Klausdorf">
          <ATHLETES>
            <ATHLETE firstname="Svantje" lastname="Glenewinkel" birthdate="2014-01-01" gender="F" nation="GER" license="448487" athleteid="34867">
              <ENTRIES>
                <ENTRY entrytime="00:12:40.15" eventid="1083" heatid="40003" lane="2">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:12:26.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.52" eventid="1123" heatid="40031" lane="6">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:33.61" />
                </ENTRY>
                <ENTRY entrytime="00:03:51.35" eventid="1163" heatid="40112" lane="1">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:03:14.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.39" eventid="1227" heatid="40197" lane="6">
                  <MEETINFO name="SHSV-Kurzbahn MS" city="Kiel" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:25.39" />
                </ENTRY>
                <ENTRY entrytime="00:06:45.95" eventid="1247" heatid="40233" lane="5">
                  <MEETINFO name="Neptun Schwimmfest" city="Kiel" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:06:45.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.56" eventid="1267" heatid="40267" lane="2">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:01:12.88" />
                </ENTRY>
                <ENTRY entrytime="00:03:26.30" eventid="1307" heatid="40348" lane="4">
                  <MEETINFO name="Bille Cup" city="Lübeck" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:03:26.30" />
                </ENTRY>
                <ENTRY entrytime="00:03:06.97" eventid="1347" heatid="40404" lane="3">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:02:50.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.59" eventid="1367" heatid="40443" lane="5">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:39.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3593" nation="GER" region="13" clubid="37045" name="SV Halle / Saale">
          <ATHLETES>
            <ATHLETE firstname="Leandro" lastname="Hanf" birthdate="2013-01-01" gender="M" nation="GER" license="464263" athleteid="37185">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.50" eventid="1133" heatid="40065" lane="3">
                  <MEETINFO name="Kids-Cup Teil 1 des LSVSA der Leistungsstützpunkte" city="Bitterfeld-Wolfen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:33.07" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.79" eventid="1173" heatid="40134" lane="3">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:49.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.53" eventid="1217" heatid="40176" lane="6">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:45.53" />
                </ENTRY>
                <ENTRY entrytime="00:05:28.58" eventid="1257" heatid="40249" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:05:28.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.31" eventid="1277" heatid="40294" lane="2">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:09.30" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.69" eventid="1317" heatid="40365" lane="7">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:59.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Tom" lastname="Kiessler" birthdate="2014-01-01" gender="M" nation="GER" license="466999" athleteid="37204">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.52" eventid="1133" heatid="40064" lane="8">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:34.52" />
                </ENTRY>
                <ENTRY entrytime="00:03:19.82" eventid="1173" heatid="40128" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:19.82" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.13" eventid="1217" heatid="40176" lane="8">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:44.68" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.00" eventid="1237" heatid="40215" lane="4">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:27.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.22" eventid="1277" heatid="40288" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:01:22.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.47" eventid="1297" heatid="40331" lane="5">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:40.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Schwenke" birthdate="2015-01-01" gender="F" nation="GER" license="450492" athleteid="37237">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.56" eventid="1123" heatid="40033" lane="5">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:33.56" />
                </ENTRY>
                <ENTRY entrytime="00:03:30.00" eventid="1163" heatid="40112" lane="2" />
                <ENTRY entrytime="00:00:41.50" eventid="1207" heatid="40164" lane="8">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:40.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.84" eventid="1267" heatid="40264" lane="8">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:01:19.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.10" eventid="1287" heatid="40314" lane="8">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:38.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.16" eventid="1327" heatid="40381" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:01:32.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Vincent" lastname="Götze" birthdate="2013-01-01" gender="M" nation="GER" license="448825" athleteid="37179">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.52" eventid="1133" heatid="40068" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:32.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.57" eventid="1173" heatid="40133" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:52.57" />
                </ENTRY>
                <ENTRY entrytime="00:05:18.98" eventid="1257" heatid="40251" lane="4">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:05:18.98" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.81" eventid="1277" heatid="40295" lane="3">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:06.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.39" eventid="1317" heatid="40368" lane="7">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:49.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emil-Friedrich" lastname="Pöpperl" birthdate="2014-01-01" gender="M" nation="GER" license="450469" athleteid="37217">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.36" eventid="1133" heatid="40062" lane="5">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:35.36" />
                </ENTRY>
                <ENTRY entrytime="00:03:14.13" eventid="1173" heatid="40129" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:14.13" />
                </ENTRY>
                <ENTRY entrytime="00:05:53.12" eventid="1257" heatid="40247" lane="3">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:05:53.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.79" eventid="1277" heatid="40290" lane="3">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:01:18.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.53" eventid="1297" heatid="40333" lane="8">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:38.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Vinz" birthdate="2013-01-01" gender="M" nation="GER" license="450459" athleteid="37244">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.95" eventid="1133" heatid="40073" lane="1">
                  <MEETINFO name="Kids-Cup Teil 1 des LSVSA der Leistungsstützpunkte" city="Bitterfeld-Wolfen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:28.65" />
                </ENTRY>
                <ENTRY entrytime="00:03:06.97" eventid="1153" heatid="40105" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:06.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.47" eventid="1217" heatid="40181" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:38.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.60" eventid="1237" heatid="40225" lane="6">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:13.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.04" eventid="1277" heatid="40302" lane="7">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:00.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.19" eventid="1297" heatid="40334" lane="8">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:30.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Jäger" birthdate="2014-01-01" gender="M" nation="GER" license="450452" athleteid="37197">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.15" eventid="1133" heatid="40066" lane="3">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:33.15" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.93" eventid="1173" heatid="40130" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:03.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.23" eventid="1237" heatid="40218" lane="7">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:24.54" />
                </ENTRY>
                <ENTRY entrytime="00:05:42.80" eventid="1257" heatid="40248" lane="7">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:05:42.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.24" eventid="1277" heatid="40293" lane="6">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:12.38" />
                </ENTRY>
                <ENTRY entrytime="00:03:11.69" eventid="1317" heatid="40363" lane="4">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:03:11.69" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Mojzis" birthdate="2015-01-01" gender="F" nation="GER" license="485022" athleteid="37211">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.74" eventid="1123" heatid="40030" lane="6">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:34.74" />
                </ENTRY>
                <ENTRY entrytime="00:03:23.79" eventid="1143" heatid="40092" lane="2">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:03:23.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.09" eventid="1207" heatid="40168" lane="4">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:37.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.30" eventid="1287" heatid="40312" lane="7">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:42.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.05" eventid="1327" heatid="40381" lane="4">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:26.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lucia Sophie" lastname="Schröter" birthdate="2013-01-01" gender="F" nation="GER" license="440281" athleteid="37230">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.55" eventid="1123" heatid="40031" lane="7">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:34.55" />
                </ENTRY>
                <ENTRY entrytime="00:03:02.45" eventid="1163" heatid="40115" lane="4">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:03:02.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.71" eventid="1227" heatid="40199" lane="2">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:21.94" />
                </ENTRY>
                <ENTRY entrytime="00:05:33.70" eventid="1247" heatid="40237" lane="3">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:05:33.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.33" eventid="1267" heatid="40266" lane="1">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:10.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.52" eventid="1307" heatid="40354" lane="5">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:53.52" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Birke" birthdate="2015-01-01" gender="F" nation="GER" license="450486" athleteid="37172">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.01" eventid="1123" heatid="40030" lane="8">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:35.01" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.88" eventid="1163" heatid="40116" lane="8">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:01.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.50" eventid="1227" heatid="40193" lane="1">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:21.77" />
                </ENTRY>
                <ENTRY entrytime="00:05:47.49" eventid="1247" heatid="40236" lane="8">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:05:47.49" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.87" eventid="1267" heatid="40266" lane="8">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:13.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.23" eventid="1287" heatid="40313" lane="4">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:37.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Elias" lastname="Quickert" birthdate="2014-01-01" gender="M" nation="GER" license="467018" athleteid="37223">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.97" eventid="1133" heatid="40063" lane="7">
                  <MEETINFO name="Kids-Cup Teil 1 des LSVSA der Leistungsstützpunkte" city="Bitterfeld-Wolfen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:33.96" />
                </ENTRY>
                <ENTRY entrytime="00:03:32.81" eventid="1153" heatid="40102" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:32.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.63" eventid="1217" heatid="40177" lane="7">
                  <MEETINFO name="1. Adventschwimmen des SV Halle" city="Halle (Saale)" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:44.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:46.78" eventid="1237" heatid="40214" lane="3">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:26.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.05" eventid="1277" heatid="40291" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-05" qualificationtime="00:01:17.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:44.06" eventid="1337" heatid="40391" lane="4">
                  <MEETINFO name="16. KBM S-A  Jg. 2012 - 2015" city="Dessau" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:36.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fiona Sophie" lastname="Hilbich" birthdate="2010-01-01" gender="F" nation="GER" license="419502" athleteid="37192">
              <ENTRIES>
                <ENTRY entrytime="00:02:42.89" eventid="1143" heatid="40099" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:42.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.62" eventid="1227" heatid="40212" lane="8">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:01:10.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.13" eventid="1287" heatid="40327" lane="5">
                  <MEETINFO name="Überprüfungswettkampf" city="Halle (Saale)" course="LCM" approved="GER" date="2025-02-08" qualificationtime="00:00:31.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.64" eventid="1327" heatid="40390" lane="5">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:01:16.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6466" nation="GER" region="12" clubid="37251" name="SSG Leipzig e.V.">
          <ATHLETES>
            <ATHLETE firstname="Emma" lastname="Zelle" birthdate="2013-01-01" gender="F" nation="GER" license="449530" athleteid="37613">
              <ENTRIES>
                <ENTRY entrytime="00:12:21.95" eventid="1083" heatid="40003" lane="6">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:12:21.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.99" eventid="1123" heatid="40040" lane="8">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:33.34" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.23" eventid="1163" heatid="40117" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:55.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.27" eventid="1227" heatid="40201" lane="1">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:01:22.27" />
                </ENTRY>
                <ENTRY entrytime="00:05:49.03" eventid="1247" heatid="40235" lane="4">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:05:49.03" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.40" eventid="1307" heatid="40355" lane="7">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:52.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:42.97" eventid="1327" heatid="40379" lane="8">
                  <MEETINFO name="Messesprintpokal des Postschwimmverein Leipzig e.V" city="Leipzig" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:01:42.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.72" eventid="1347" heatid="40408" lane="1">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:44.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.26" eventid="1387" heatid="40481" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:17.26" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nele" lastname="Clauß" birthdate="2008-01-01" gender="F" nation="GER" license="366218" athleteid="37304">
              <ENTRIES>
                <ENTRY entrytime="00:05:19.64" eventid="1063" heatid="39997" lane="1">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-14" qualificationtime="00:05:19.64" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.21" eventid="1143" heatid="40097" lane="2" />
                <ENTRY entrytime="00:00:38.95" eventid="1207" heatid="40169" lane="8">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:39.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.01" eventid="1227" heatid="40210" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marlon" lastname="Jung" birthdate="2009-01-01" gender="M" nation="GER" license="391282" athleteid="37375">
              <HANDICAP exception="12+" />
              <ENTRIES>
                <ENTRY entrytime="00:09:23.35" eventid="1093" heatid="40018" lane="3">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:09:23.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.64" eventid="1133" heatid="40077" lane="8" />
                <ENTRY entrytime="00:02:41.08" eventid="1173" heatid="40136" lane="5" />
                <ENTRY entrytime="00:02:26.06" eventid="1197" heatid="40155" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:26.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.37" eventid="1217" heatid="40186" lane="2">
                  <MEETINFO name="DKM Para Schwimmen offen für DSV-Schwimmer" city="Nürnberg" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:00:34.37" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.58" eventid="1277" heatid="40306" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:59.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.94" eventid="1317" heatid="40375" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:21.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.14" eventid="1397" heatid="40495" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:04.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Phoebe" lastname="Lißner" birthdate="2013-01-01" gender="F" nation="GER" license="448337" athleteid="37425">
              <ENTRIES>
                <ENTRY entrytime="00:10:46.94" eventid="1083" heatid="40008" lane="5" />
                <ENTRY entrytime="00:00:31.70" eventid="1123" heatid="40042" lane="5" />
                <ENTRY entrytime="00:03:00.25" eventid="1143" heatid="40097" lane="3">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:00.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.57" eventid="1207" heatid="40161" lane="1" />
                <ENTRY entrytime="00:04:55.16" eventid="1247" heatid="40243" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:04:55.16" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.39" eventid="1287" heatid="40327" lane="7">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:31.39" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.62" eventid="1327" heatid="40389" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:01:27.11" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.03" eventid="1347" heatid="40418" lane="8">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:21.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.67" eventid="1367" heatid="40456" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:33.67" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alexander" lastname="Belyavskiy" birthdate="2010-01-01" gender="M" nation="GER" license="426136" athleteid="37260">
              <ENTRIES>
                <ENTRY entrytime="00:17:37.94" eventid="1113" heatid="40025" lane="5" />
                <ENTRY entrytime="00:03:06.19" eventid="1153" heatid="40105" lane="4" />
                <ENTRY entrytime="00:02:18.17" eventid="1197" heatid="40156" lane="7">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:02:18.17" />
                </ENTRY>
                <ENTRY entrytime="00:04:26.47" eventid="1257" heatid="40259" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:04:26.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.47" eventid="1277" heatid="40306" lane="4">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:59.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.06" eventid="1317" heatid="40375" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:20.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.25" eventid="1357" heatid="40437" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:02.25" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.03" eventid="1397" heatid="40496" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:01.96" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Wießner" birthdate="2012-01-01" gender="F" nation="GER" license="434536" athleteid="37603">
              <ENTRIES>
                <ENTRY entrytime="00:11:01.31" eventid="1083" heatid="40007" lane="7" />
                <ENTRY entrytime="00:00:27.93" eventid="1123" heatid="40057" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.93" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.13" eventid="1163" heatid="40122" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:43.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.29" eventid="1207" heatid="40168" lane="8">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:00:39.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.69" eventid="1227" heatid="40210" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:15.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.00" eventid="1307" heatid="40358" lane="7">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:41.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.47" eventid="1327" heatid="40383" lane="4">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:01:31.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.10" eventid="1367" heatid="40457" lane="7">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:33.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.26" eventid="1387" heatid="40484" lane="6">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:01:15.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Frederik Alexander" lastname="Kaul" birthdate="2011-01-01" gender="M" nation="GER" license="416013" athleteid="37384">
              <ENTRIES>
                <ENTRY entrytime="00:09:12.74" eventid="1093" heatid="40018" lane="5">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:09:12.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.52" eventid="1133" heatid="40074" lane="4">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:29.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.92" eventid="1153" heatid="40107" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:55.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.37" eventid="1217" heatid="40179" lane="6">
                  <MEETINFO name="Jugend trainiert für Olympia - Sachsen" city="Leipzig" course="LCM" approved="GER" date="2025-03-20" qualificationtime="00:00:40.37" />
                </ENTRY>
                <ENTRY entrytime="00:04:31.93" eventid="1257" heatid="40258" lane="5">
                  <MEETINFO name="17. Helfmann-Cup" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:04:26.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.32" eventid="1277" heatid="40305" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:00.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.06" eventid="1317" heatid="40373" lane="7">
                  <MEETINFO name="17. Helfmann-Cup" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:02:26.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.93" eventid="1357" heatid="40436" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:07.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.39" eventid="1377" heatid="40470" lane="1">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:33.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Severyuk" birthdate="2012-01-01" gender="M" nation="GER" license="440973" athleteid="37545">
              <ENTRIES>
                <ENTRY entrytime="00:05:42.95" eventid="1073" heatid="40000" lane="1" />
                <ENTRY entrytime="00:00:27.27" eventid="1133" heatid="40081" lane="4">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:28.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.25" eventid="1173" heatid="40141" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:19.25" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.19" eventid="1197" heatid="40152" lane="5" />
                <ENTRY entrytime="00:04:58.39" eventid="1257" heatid="40255" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:04:58.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.81" eventid="1277" heatid="40308" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:58.98" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.05" eventid="1337" heatid="40395" lane="7">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:01:32.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.26" eventid="1357" heatid="40435" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:10.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.25" eventid="1397" heatid="40495" lane="8">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:01:05.22" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fabian" lastname="Brauer" birthdate="2013-01-01" gender="M" nation="GER" license="445392" athleteid="37284">
              <ENTRIES>
                <ENTRY entrytime="00:10:37.67" eventid="1093" heatid="40015" lane="1" />
                <ENTRY entrytime="00:00:27.97" eventid="1133" heatid="40079" lane="3">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:27.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.76" eventid="1173" heatid="40138" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:35.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.50" eventid="1197" heatid="40154" lane="6">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:33.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.49" eventid="1237" heatid="40227" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:01:12.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.12" eventid="1297" heatid="40341" lane="6">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:30.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.38" eventid="1337" heatid="40399" lane="6">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:22.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.57" eventid="1377" heatid="40469" lane="3">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:33.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.04" eventid="1397" heatid="40493" lane="7">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:08.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Niklas" lastname="Turich" birthdate="2010-01-01" gender="M" nation="GER" license="417679" athleteid="37584">
              <ENTRIES>
                <ENTRY entrytime="00:05:53.80" eventid="1073" heatid="39999" lane="6" />
                <ENTRY entrytime="00:02:39.89" eventid="1153" heatid="40110" lane="7">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:02:39.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.49" eventid="1197" heatid="40152" lane="3" />
                <ENTRY entrytime="00:04:35.88" eventid="1257" heatid="40258" lane="6">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:04:43.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.82" eventid="1277" heatid="40304" lane="3" />
                <ENTRY entrytime="00:01:11.19" eventid="1337" heatid="40402" lane="7">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-25" qualificationtime="00:01:11.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.01" eventid="1357" heatid="40434" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:12.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.59" eventid="1397" heatid="40494" lane="3">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:04.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Harnisch" birthdate="2010-01-01" gender="M" nation="GER" license="406011" athleteid="37332">
              <ENTRIES>
                <ENTRY entrytime="00:04:56.09" eventid="1073" heatid="40001" lane="3">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:04:57.61" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.49" eventid="1133" heatid="40087" lane="7">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:26.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.49" eventid="1197" heatid="40154" lane="3" />
                <ENTRY entrytime="00:04:16.70" eventid="1257" heatid="40259" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:04:16.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.00" eventid="1277" heatid="40311" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:55.25" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.32" eventid="1317" heatid="40375" lane="5">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:02:20.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.51" eventid="1357" heatid="40438" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:01.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Aaliyah" lastname="Schiffel" birthdate="2006-01-01" gender="F" nation="GER" license="348758" athleteid="37495">
              <ENTRIES>
                <ENTRY entrytime="00:09:29.11" eventid="1083" heatid="40011" lane="3">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:09:30.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.18" eventid="1123" heatid="40056" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.04" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.92" eventid="1163" heatid="40127" lane="5" />
                <ENTRY entrytime="00:00:33.64" eventid="1207" heatid="40173" lane="4">
                  <MEETINFO name="136. Deutsche Meisterschaften im Schwimmen" city="Berlin" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:34.04" />
                </ENTRY>
                <ENTRY entrytime="00:04:42.40" eventid="1247" heatid="40245" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Malin" lastname="Petzold" birthdate="2013-01-01" gender="F" nation="GER" license="445609" athleteid="37470">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.72" eventid="1123" heatid="40042" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:31.65" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.54" eventid="1143" heatid="40096" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:03:01.25" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.92" eventid="1227" heatid="40195" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:29.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.02" eventid="1287" heatid="40316" lane="6">
                  <MEETINFO name="Plauener Herbst- Mehrkampf" city="Plauen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:34.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.45" eventid="1327" heatid="40387" lane="4">
                  <MEETINFO name="Plauener Herbst- Mehrkampf" city="Plauen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:22.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.77" eventid="1387" heatid="40480" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:01:18.77" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Leonhardt" birthdate="2014-01-01" gender="F" nation="GER" license="446794" athleteid="37407">
              <ENTRIES>
                <ENTRY entrytime="00:11:01.48" eventid="1083" heatid="40007" lane="1">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:11:01.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.24" eventid="1123" heatid="40054" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:29.24" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.66" eventid="1163" heatid="40126" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:32.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.93" eventid="1207" heatid="40173" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:34.93" />
                </ENTRY>
                <ENTRY entrytime="00:05:00.10" eventid="1247" heatid="40242" lane="4">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:00.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.10" eventid="1267" heatid="40283" lane="2">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:02.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.60" eventid="1307" heatid="40360" lane="4">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:30.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.74" eventid="1367" heatid="40456" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:33.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.25" eventid="1387" heatid="40484" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:11.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jasper" lastname="Müller" birthdate="2013-01-01" gender="M" nation="GER" license="441004" athleteid="37460">
              <ENTRIES>
                <ENTRY entrytime="00:06:32.56" eventid="1073" heatid="39998" lane="7" />
                <ENTRY entrytime="00:00:31.64" eventid="1133" heatid="40069" lane="4">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:31.64" />
                </ENTRY>
                <ENTRY entrytime="00:03:10.81" eventid="1153" heatid="40105" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:03:10.81" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.17" eventid="1197" heatid="40153" lane="7" />
                <ENTRY entrytime="00:00:42.44" eventid="1217" heatid="40178" lane="3">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:42.60" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.51" eventid="1317" heatid="40371" lane="5">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-08" qualificationtime="00:02:36.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.79" eventid="1337" heatid="40396" lane="6" />
                <ENTRY entrytime="00:00:33.88" eventid="1377" heatid="40469" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:33.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.42" eventid="1397" heatid="40491" lane="2">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:15.19" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hannah Grete" lastname="Hunger" birthdate="2013-01-01" gender="F" nation="GER" license="453218" athleteid="37365">
              <ENTRIES>
                <ENTRY entrytime="00:06:11.84" eventid="1063" heatid="39994" lane="2">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-14" qualificationtime="00:06:11.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.89" eventid="1123" heatid="40041" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:33.66" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.33" eventid="1143" heatid="40096" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:03:03.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.28" eventid="1207" heatid="40168" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:39.28" />
                </ENTRY>
                <ENTRY entrytime="00:05:22.80" eventid="1247" heatid="40238" lane="3">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:22.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.49" eventid="1267" heatid="40272" lane="2">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:10.49" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.01" eventid="1307" heatid="40356" lane="5">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:02:48.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.56" eventid="1367" heatid="40442" lane="6">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:40.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.48" eventid="1387" heatid="40479" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:20.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emma" lastname="Färber" birthdate="2011-01-01" gender="F" nation="GER" license="408425" athleteid="37314">
              <ENTRIES>
                <ENTRY entrytime="00:05:07.85" eventid="1063" heatid="39997" lane="5">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:05:07.85" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.65" eventid="1143" heatid="40099" lane="3">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:42.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.59" eventid="1207" heatid="40172" lane="6">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:36.59" />
                </ENTRY>
                <ENTRY entrytime="00:04:51.25" eventid="1247" heatid="40244" lane="7" />
                <ENTRY entrytime="00:01:01.53" eventid="1267" heatid="40285" lane="7">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:01:04.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.39" eventid="1307" heatid="40361" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:25.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.71" eventid="1347" heatid="40418" lane="7" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Janek Thorben" lastname="Reyher" birthdate="2007-01-01" gender="M" nation="GER" license="361329" athleteid="37477">
              <ENTRIES>
                <ENTRY entrytime="00:04:29.93" eventid="1073" heatid="40002" lane="4">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:04:19.74" />
                </ENTRY>
                <ENTRY entrytime="00:16:01.44" eventid="1113" heatid="40025" lane="4">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-25" qualificationtime="00:16:01.44" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.98" eventid="1173" heatid="40142" lane="3" />
                <ENTRY entrytime="00:04:06.02" eventid="1257" heatid="40260" lane="4">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:04:06.02" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.51" eventid="1317" heatid="40376" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:06.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:59.03" eventid="1357" heatid="40438" lane="3">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:59.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.91" eventid="1377" heatid="40474" lane="2">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-25" qualificationtime="00:00:27.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mara" lastname="Hacker" birthdate="2012-01-01" gender="F" nation="GER" license="440971" athleteid="37322">
              <ENTRIES>
                <ENTRY entrytime="00:11:25.22" eventid="1083" heatid="40005" lane="4">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:11:25.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.44" eventid="1123" heatid="40048" lane="3">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:00:30.44" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.79" eventid="1163" heatid="40120" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:49.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.18" eventid="1207" heatid="40168" lane="3">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:39.18" />
                </ENTRY>
                <ENTRY entrytime="00:05:24.40" eventid="1247" heatid="40238" lane="6">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:05:24.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.41" eventid="1267" heatid="40280" lane="5">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:01:07.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.07" eventid="1327" heatid="40382" lane="5">
                  <MEETINFO name="Messesprintpokal des Postschwimmverein Leipzig e.V" city="Leipzig" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:01:31.07" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.37" eventid="1347" heatid="40414" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:29.37" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.51" eventid="1387" heatid="40483" lane="1">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:13.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Justus Georg" lastname="Schüller" birthdate="2010-01-01" gender="M" nation="GER" license="396360" athleteid="37535">
              <ENTRIES>
                <ENTRY entrytime="00:09:03.70" eventid="1093" heatid="40019" lane="8">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:09:29.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.09" eventid="1133" heatid="40087" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:25.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.79" eventid="1173" heatid="40141" lane="5" />
                <ENTRY entrytime="00:02:21.03" eventid="1197" heatid="40155" lane="6">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:02:21.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.06" eventid="1217" heatid="40181" lane="5" />
                <ENTRY entrytime="00:04:14.48" eventid="1257" heatid="40260" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:04:14.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.32" eventid="1277" heatid="40310" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:55.87" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.31" eventid="1317" heatid="40373" lane="6" />
                <ENTRY entrytime="00:02:00.53" eventid="1357" heatid="40438" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:00.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jonas" lastname="Lehmann" birthdate="2014-01-01" gender="M" nation="GER" license="449099" athleteid="37404">
              <ENTRIES>
                <ENTRY entrytime="00:12:25.03" eventid="1093" heatid="40012" lane="3" />
                <ENTRY entrytime="00:05:27.48" eventid="1257" heatid="40250" lane="7">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:27.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lius Pepe" lastname="Baumeister" birthdate="2009-01-01" gender="M" nation="GER" license="391171" athleteid="37252">
              <ENTRIES>
                <ENTRY entrytime="00:04:37.26" eventid="1073" heatid="40002" lane="3">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:04:27.66" />
                </ENTRY>
                <ENTRY entrytime="00:08:25.59" eventid="1093" heatid="40019" lane="4" />
                <ENTRY entrytime="00:02:18.20" eventid="1153" heatid="40111" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:18.20" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.36" eventid="1173" heatid="40142" lane="2">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:12.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.21" eventid="1217" heatid="40190" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:29.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.44" eventid="1237" heatid="40232" lane="7">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:00:59.85" />
                </ENTRY>
                <ENTRY entrytime="00:04:07.00" eventid="1257" heatid="40260" lane="5">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:04:09.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jonas" lastname="Herrmann" birthdate="2007-01-01" gender="M" nation="GER" license="366274" athleteid="37350">
              <ENTRIES>
                <ENTRY entrytime="00:08:38.92" eventid="1093" heatid="40019" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:08:16.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.22" eventid="1133" heatid="40085" lane="7">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:26.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.67" eventid="1173" heatid="40142" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:14.67" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.33" eventid="1237" heatid="40231" lane="2">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:01:03.33" />
                </ENTRY>
                <ENTRY entrytime="00:04:12.53" eventid="1257" heatid="40260" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:04:03.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Finn" lastname="Schoop" birthdate="2011-01-01" gender="M" nation="GER" license="419064" athleteid="37521">
              <ENTRIES>
                <ENTRY entrytime="00:05:08.43" eventid="1073" heatid="40001" lane="7">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:05:08.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.03" eventid="1133" heatid="40086" lane="8">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:26.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.44" eventid="1173" heatid="40142" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:14.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.57" eventid="1237" heatid="40231" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:01.57" />
                </ENTRY>
                <ENTRY entrytime="00:04:42.48" eventid="1257" heatid="40257" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:04:42.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.40" eventid="1277" heatid="40309" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:57.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.42" eventid="1317" heatid="40376" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:17.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.38" eventid="1397" heatid="40494" lane="4">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:04.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Louis" lastname="Schubert" birthdate="2004-01-01" gender="M" nation="GER" license="358844" athleteid="37530">
              <ENTRIES>
                <ENTRY entrytime="00:04:45.09" eventid="1073" heatid="40002" lane="2" />
                <ENTRY entrytime="00:00:22.86" eventid="1133" heatid="40089" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:23.47" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.64" eventid="1153" heatid="40110" lane="8" />
                <ENTRY entrytime="NT" eventid="1237" heatid="40214" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Carlotta" lastname="Waizmann" birthdate="2009-01-01" gender="F" nation="GER" license="391769" athleteid="37593">
              <ENTRIES>
                <ENTRY entrytime="00:09:35.04" eventid="1083" heatid="40011" lane="6">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:09:37.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.32" eventid="1123" heatid="40058" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.14" eventid="1163" heatid="40126" lane="5" />
                <ENTRY entrytime="00:02:15.66" eventid="1187" heatid="40150" lane="4">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-13" qualificationtime="00:02:15.66" />
                </ENTRY>
                <ENTRY entrytime="00:04:40.69" eventid="1247" heatid="40245" lane="7" />
                <ENTRY entrytime="00:00:28.04" eventid="1287" heatid="40329" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:28.28" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.56" eventid="1307" heatid="40361" lane="4">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:20.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.91" eventid="1347" heatid="40420" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:06.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.51" eventid="1387" heatid="40485" lane="4">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:01:01.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mads Jakob" lastname="Strauch" birthdate="2013-01-01" gender="M" nation="GER" license="445296" athleteid="37564">
              <ENTRIES>
                <ENTRY entrytime="00:11:18.71" eventid="1093" heatid="40013" lane="1" />
                <ENTRY entrytime="00:00:32.40" eventid="1133" heatid="40068" lane="7">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:32.40" />
                </ENTRY>
                <ENTRY entrytime="00:03:12.00" eventid="1153" heatid="40104" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:12.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.16" eventid="1217" heatid="40176" lane="4">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:45.16" />
                </ENTRY>
                <ENTRY entrytime="00:05:02.31" eventid="1257" heatid="40254" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:05:02.31" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.89" eventid="1317" heatid="40368" lane="5">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-08" qualificationtime="00:02:47.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.97" eventid="1337" heatid="40395" lane="5">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:29.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.54" eventid="1357" heatid="40429" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:24.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.31" eventid="1397" heatid="40488" lane="3">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:25.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mercedesz" lastname="Lißner" birthdate="2010-01-01" gender="F" nation="GER" license="426137" athleteid="37417">
              <ENTRIES>
                <ENTRY entrytime="00:10:06.09" eventid="1083" heatid="40010" lane="6">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:10:06.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.30" eventid="1123" heatid="40056" lane="7">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:28.96" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.59" eventid="1163" heatid="40127" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:23.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.30" eventid="1227" heatid="40213" lane="5" />
                <ENTRY entrytime="00:00:59.96" eventid="1267" heatid="40286" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:00.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.89" eventid="1307" heatid="40361" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:25.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.53" eventid="1347" heatid="40420" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:10.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Florin" lastname="Thomas" birthdate="2013-01-01" gender="M" nation="GER" license="437788" athleteid="37574">
              <ENTRIES>
                <ENTRY entrytime="00:11:37.32" eventid="1093" heatid="40013" lane="8" />
                <ENTRY entrytime="00:00:30.62" eventid="1133" heatid="40071" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:00:30.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.05" eventid="1173" heatid="40136" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:42.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.60" eventid="1197" heatid="40152" lane="7">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:02:58.60" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.01" eventid="1237" heatid="40222" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:01:20.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.01" eventid="1277" heatid="40301" lane="8">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:05.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.67" eventid="1317" heatid="40372" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:35.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.22" eventid="1377" heatid="40465" lane="1">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:37.22" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.14" eventid="1397" heatid="40490" lane="7">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:17.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anna Franziska" lastname="Hunger" birthdate="2011-01-01" gender="F" nation="GER" license="428578" athleteid="37356">
              <ENTRIES>
                <ENTRY entrytime="00:05:08.34" eventid="1063" heatid="39997" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:05:08.34" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.22" eventid="1143" heatid="40099" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:39.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.54" eventid="1207" heatid="40173" lane="2">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:36.08" />
                </ENTRY>
                <ENTRY entrytime="00:04:53.27" eventid="1247" heatid="40244" lane="8">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:04:53.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.63" eventid="1267" heatid="40286" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:00.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.68" eventid="1307" heatid="40361" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:24.68" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.62" eventid="1347" heatid="40416" lane="5" />
                <ENTRY entrytime="00:00:33.47" eventid="1367" heatid="40457" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Carl" lastname="Brückner" birthdate="2014-01-01" gender="M" nation="GER" license="454910" athleteid="37294">
              <ENTRIES>
                <ENTRY entrytime="00:12:08.11" eventid="1093" heatid="40012" lane="5" />
                <ENTRY entrytime="00:00:31.48" eventid="1133" heatid="40070" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:32.17" />
                </ENTRY>
                <ENTRY entrytime="00:03:27.80" eventid="1153" heatid="40103" lane="7">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:03:27.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.83" eventid="1217" heatid="40176" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:45.83" />
                </ENTRY>
                <ENTRY entrytime="00:05:17.57" eventid="1257" heatid="40252" lane="1">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:17.57" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.65" eventid="1317" heatid="40369" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:47.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.62" eventid="1337" heatid="40394" lane="2">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:33.62" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.14" eventid="1357" heatid="40427" lane="7">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:33.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.63" eventid="1377" heatid="40465" lane="8">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:37.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Möschke" birthdate="2013-01-01" gender="F" nation="GER" license="448338" athleteid="37450">
              <ENTRIES>
                <ENTRY entrytime="00:11:13.99" eventid="1083" heatid="40006" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:11:13.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.92" eventid="1123" heatid="40040" lane="6">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:00:31.92" />
                </ENTRY>
                <ENTRY entrytime="00:03:16.88" eventid="1143" heatid="40093" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:16.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.89" eventid="1207" heatid="40161" lane="3">
                  <MEETINFO name="Jugend trainiert für Olympia - Sachsen" city="Leipzig" course="LCM" approved="GER" date="2025-03-20" qualificationtime="00:00:41.47" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.53" eventid="1227" heatid="40207" lane="4">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:01:16.14" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.15" eventid="1267" heatid="40275" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:10.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.12" eventid="1327" heatid="40384" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:01:36.01" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.37" eventid="1347" heatid="40412" lane="5">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:33.37" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.24" eventid="1367" heatid="40455" lane="1">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:34.24" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Rosa" lastname="Schindler" birthdate="2012-01-01" gender="F" nation="GER" license="440950" athleteid="37501">
              <ENTRIES>
                <ENTRY entrytime="00:10:37.78" eventid="1083" heatid="40009" lane="6">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:10:37.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.55" eventid="1123" heatid="40043" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:31.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.31" eventid="1163" heatid="40120" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:48.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.95" eventid="1207" heatid="40158" lane="5" />
                <ENTRY entrytime="00:01:18.36" eventid="1227" heatid="40204" lane="5">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:01:18.36" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.63" eventid="1267" heatid="40273" lane="4">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:01:09.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.08" eventid="1307" heatid="40356" lane="2">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:49.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.52" eventid="1367" heatid="40452" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:35.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.56" eventid="1387" heatid="40481" lane="4">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:01:15.56" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Frida" lastname="Meißner" birthdate="2014-01-01" gender="F" nation="GER" license="448123" athleteid="37440">
              <ENTRIES>
                <ENTRY entrytime="00:11:28.95" eventid="1083" heatid="40005" lane="2">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:11:28.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.04" eventid="1123" heatid="40050" lane="1">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:00:31.45" />
                </ENTRY>
                <ENTRY entrytime="00:03:19.50" eventid="1143" heatid="40092" lane="4">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:19.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.77" eventid="1207" heatid="40160" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:44.78" />
                </ENTRY>
                <ENTRY entrytime="00:05:17.39" eventid="1247" heatid="40240" lane="1">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:17.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.12" eventid="1287" heatid="40322" lane="5">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:32.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.05" eventid="1327" heatid="40381" lane="7">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:34.05" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.69" eventid="1367" heatid="40451" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:35.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.25" eventid="1387" heatid="40482" lane="2">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:15.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Luschnitz" birthdate="2008-01-01" gender="F" nation="GER" license="389677" athleteid="37435">
              <ENTRIES>
                <ENTRY entrytime="00:09:35.14" eventid="1083" heatid="40011" lane="2">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:09:35.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.78" eventid="1123" heatid="40058" lane="6" />
                <ENTRY entrytime="00:02:26.68" eventid="1163" heatid="40127" lane="2" />
                <ENTRY entrytime="00:01:06.34" eventid="1227" heatid="40213" lane="3">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:05.09" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Helena Sophie" lastname="Haupt" birthdate="2012-01-01" gender="F" nation="GER" license="443234" athleteid="37340">
              <ENTRIES>
                <ENTRY entrytime="00:05:43.06" eventid="1063" heatid="39996" lane="3">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-14" qualificationtime="00:05:43.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.97" eventid="1123" heatid="40055" lane="1">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:28.97" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.67" eventid="1143" heatid="40096" lane="6">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:03:03.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.78" eventid="1207" heatid="40171" lane="8">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:37.78" />
                </ENTRY>
                <ENTRY entrytime="00:05:11.92" eventid="1247" heatid="40241" lane="4">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:05:11.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.63" eventid="1267" heatid="40285" lane="8">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:01:03.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.21" eventid="1307" heatid="40359" lane="6">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:36.21" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.84" eventid="1347" heatid="40417" lane="3">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:22.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.05" eventid="1387" heatid="40480" lane="2">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:01:18.24" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mick Günter" lastname="Birgel" birthdate="2012-01-01" gender="M" nation="GER" license="407310" athleteid="37269">
              <ENTRIES>
                <ENTRY entrytime="00:11:45.12" eventid="1093" heatid="40012" lane="4" />
                <ENTRY entrytime="00:00:26.85" eventid="1133" heatid="40084" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:26.85" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.69" eventid="1153" heatid="40108" lane="7">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:52.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.10" eventid="1217" heatid="40182" lane="4">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:37.44" />
                </ENTRY>
                <ENTRY entrytime="00:04:45.00" eventid="1257" heatid="40256" lane="2">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:04:45.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.13" eventid="1297" heatid="40344" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:28.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.05" eventid="1337" heatid="40401" lane="6">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:22.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.52" eventid="1357" heatid="40434" lane="2">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:12.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.46" eventid="1397" heatid="40495" lane="2">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:01:01.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ronja" lastname="Stodolka" birthdate="2010-01-01" gender="F" nation="GER" license="406010" athleteid="37555">
              <ENTRIES>
                <ENTRY entrytime="00:10:27.16" eventid="1083" heatid="40009" lane="5">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:10:27.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.20" eventid="1143" heatid="40099" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:42.20" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.34" eventid="1187" heatid="40150" lane="6" />
                <ENTRY entrytime="00:01:10.89" eventid="1227" heatid="40211" lane="5">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:01:13.31" />
                </ENTRY>
                <ENTRY entrytime="00:05:15.51" eventid="1247" heatid="40240" lane="6" />
                <ENTRY entrytime="00:02:26.29" eventid="1307" heatid="40361" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:27.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.48" eventid="1367" heatid="40454" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:34.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.87" eventid="1387" heatid="40485" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:09.67" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Limaris" lastname="Dix" birthdate="2007-01-01" gender="M" nation="GER" license="376786" athleteid="37309">
              <ENTRIES>
                <ENTRY entrytime="00:04:45.25" eventid="1073" heatid="40002" lane="7" />
                <ENTRY entrytime="00:00:22.70" eventid="1133" heatid="40089" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:23.36" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.91" eventid="1197" heatid="40156" lane="6">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:02:08.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.64" eventid="1217" heatid="40188" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ben" lastname="Bodusch" birthdate="2008-01-01" gender="M" nation="GER" license="377824" athleteid="37279">
              <ENTRIES>
                <ENTRY entrytime="00:04:34.18" eventid="1073" heatid="40002" lane="5">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:04:21.77" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.07" eventid="1173" heatid="40142" lane="6" />
                <ENTRY entrytime="00:00:31.07" eventid="1217" heatid="40189" lane="2">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-27" qualificationtime="00:00:31.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.58" eventid="1237" heatid="40232" lane="3">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:01:00.34" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Justus" lastname="Richter" birthdate="2013-01-01" gender="M" nation="GER" license="444299" athleteid="37485">
              <ENTRIES>
                <ENTRY entrytime="00:05:46.25" eventid="1073" status="WDR" heatid="39999" lane="4">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-14" qualificationtime="00:05:46.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.51" eventid="1133" status="WDR" heatid="40070" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:31.51" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.79" eventid="1173" status="WDR" heatid="40137" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:38.79" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.99" eventid="1197" status="WDR" heatid="40152" lane="1">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:03:00.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.27" eventid="1237" status="WDR" heatid="40224" lane="2">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:01:18.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.30" eventid="1277" status="WDR">
                  <MEETINFO name="Messesprintpokal des Postschwimmverein Leipzig e.V" city="Leipzig" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:01:09.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.23" eventid="1317" status="WDR">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:38.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.21" eventid="1377" status="WDR">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:36.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.33" eventid="1397" status="WDR">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:19.33" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Julia Franziska" lastname="Kaul" birthdate="2011-01-01" gender="F" nation="GER" license="416012" athleteid="37394">
              <ENTRIES>
                <ENTRY entrytime="00:05:14.45" eventid="1063" heatid="39997" lane="2">
                  <MEETINFO name="HM und HJM Langbahn  Darmstadt" city="Darmstadt" course="LCM" approved="GER" date="2025-06-20" qualificationtime="00:05:14.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.29" eventid="1123" heatid="40053" lane="4">
                  <MEETINFO name="Jugend trainert für Olympia" city="Berlin" course="SCM" approved="GER" date="2025-09-23" qualificationtime="00:00:28.47" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.25" eventid="1163" heatid="40126" lane="3">
                  <MEETINFO name="17. Helfmann-Cup" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:02:29.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.50" eventid="1207" heatid="40167" lane="7">
                  <MEETINFO name="Jugend trainert für Olympia" city="Berlin" course="SCM" approved="GER" date="2025-09-23" qualificationtime="00:00:40.58" />
                </ENTRY>
                <ENTRY entrytime="00:04:26.12" eventid="1247" heatid="40245" lane="3">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:04:26.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.55" eventid="1287" heatid="40329" lane="8">
                  <MEETINFO name="BaHaMa Cup" city="Langen" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:00:30.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.41" eventid="1327" heatid="40383" lane="1" />
                <ENTRY entrytime="00:00:34.98" eventid="1367" heatid="40453" lane="4">
                  <MEETINFO name="17. Helfmann-Cup" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-02-02" qualificationtime="00:00:34.17" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.62" eventid="1387" heatid="40485" lane="2">
                  <MEETINFO name="HM und HJM Langbahn  Darmstadt" city="Darmstadt" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:06.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ninett" lastname="Schönberg" birthdate="2011-01-01" gender="F" nation="GER" license="418811" athleteid="37511">
              <ENTRIES>
                <ENTRY entrytime="00:05:32.30" eventid="1063" status="WDR" heatid="39996" lane="5" />
                <ENTRY entrytime="00:00:27.38" eventid="1123" status="WDR" heatid="40058" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.38" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.97" eventid="1163" status="WDR" heatid="40124" lane="1">
                  <MEETINFO name="34. Hallescher Salzpokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-10-04" qualificationtime="00:02:39.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.32" eventid="1187" status="WDR" heatid="40149" lane="4">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:40.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.48" eventid="1227" status="WDR" heatid="40212" lane="1">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:01:14.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.58" eventid="1287" status="WDR">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:30.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.37" eventid="1327" status="WDR">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:01:20.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.53" eventid="1367" status="WDR">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:00:33.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.09" eventid="1387" status="WDR">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:10.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="37994" name="SK Motorlet Praha">
          <CONTACT email="skmop@skmop.cz" internet="www.skmop.cz" name="SK Motorlet Praha, spolek" street="Radlická 298/105" street2="Praha 5" zip="15500" />
          <ATHLETES>
            <ATHLETE firstname="Matfej" lastname="Krychfalushiy" birthdate="2013-07-13" gender="M" nation="UKR" athleteid="38025">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.30" entrycourse="SCM" eventid="1133" heatid="40068" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:53.15" entrycourse="SCM" eventid="1173" heatid="40133" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:01:21.93" entrycourse="SCM" eventid="1237" heatid="40221" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:05:31.38" entrycourse="SCM" eventid="1257" heatid="40249" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:01:12.52" entrycourse="SCM" eventid="1277" heatid="40294" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:00:42.43" entrycourse="SCM" eventid="1297" heatid="40332" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:02:42.06" entrycourse="SCM" eventid="1357" heatid="40424" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:39.03" entrycourse="SCM" eventid="1377" heatid="40464" lane="8">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Petr" lastname="Liška" birthdate="2013-01-16" gender="M" nation="CZE" athleteid="38034">
              <ENTRIES>
                <ENTRY entrytime="00:05:52.50" entrycourse="SCM" eventid="1073" heatid="39999" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:29.67" entrycourse="SCM" eventid="1133" heatid="40074" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:55.30" entrycourse="SCM" eventid="1153" heatid="40107" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:02:28.65" entrycourse="SCM" eventid="1173" heatid="40139" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:00:37.40" entrycourse="SCM" eventid="1217" heatid="40182" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:01:09.77" entrycourse="SCM" eventid="1237" heatid="40229" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:05:02.00" entrycourse="SCM" eventid="1257" heatid="40254" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:04.25" entrycourse="SCM" eventid="1277" heatid="40300" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:33.81" entrycourse="SCM" eventid="1297" heatid="40336" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:01:20.52" entrycourse="SCM" eventid="1337" heatid="40398" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:32.04" entrycourse="SCM" eventid="1377" heatid="40471" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:01:22.00" entrycourse="SCM" eventid="1397" heatid="40489" lane="8">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Gryč" birthdate="2012-10-12" gender="M" nation="CZE" athleteid="38018">
              <ENTRIES>
                <ENTRY entrytime="00:20:19.15" entrycourse="SCM" eventid="1113" heatid="40024" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:00:29.19" entrycourse="SCM" eventid="1133" heatid="40075" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:02:49.42" entrycourse="SCM" eventid="1173" heatid="40135" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:05:04.87" entrycourse="SCM" eventid="1257" heatid="40254" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:04.66" entrycourse="SCM" eventid="1277" heatid="40300" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:02:21.65" entrycourse="SCM" eventid="1357" heatid="40430" lane="5">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Julie" lastname="Zusková" birthdate="2012-04-13" gender="F" nation="CZE" athleteid="38083">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.58" entrycourse="SCM" eventid="1123" status="WDR" heatid="40048" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:02:41.29" entrycourse="SCM" eventid="1163" status="WDR" heatid="40123" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:01:14.26" entrycourse="SCM" eventid="1227" status="WDR" heatid="40209" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:01:07.52" entrycourse="SCM" eventid="1267" status="WDR">
                </ENTRY>
                <ENTRY entrytime="00:00:33.48" entrycourse="SCM" eventid="1287" status="WDR">
                </ENTRY>
                <ENTRY entrytime="00:02:42.59" entrycourse="SCM" eventid="1307" status="WDR">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Makar" lastname="Fijal" birthdate="2013-10-13" gender="M" nation="UKR" athleteid="38014">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.97" entrycourse="SCM" eventid="1277" heatid="40292" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:03:14.52" entrycourse="SCM" eventid="1317" heatid="40363" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:01:27.09" entrycourse="SCM" eventid="1397" heatid="40488" lane="2">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Matyáš Hugo" lastname="Března" birthdate="2015-12-31" gender="M" nation="CZE" athleteid="38002">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" entrycourse="SCM" eventid="1133" heatid="40059" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:00:49.00" entrycourse="SCM" eventid="1217" heatid="40174" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:01:38.10" entrycourse="SCM" eventid="1277" heatid="40287" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:01:47.14" entrycourse="SCM" eventid="1337" heatid="40391" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:48.31" entrycourse="SCM" eventid="1377" heatid="40460" lane="5">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nela" lastname="Zugarová" birthdate="2013-07-12" gender="F" nation="CZE" athleteid="38076">
              <ENTRIES>
                <ENTRY entrytime="00:11:01.16" entrycourse="SCM" eventid="1083" heatid="40007" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:31.91" entrycourse="SCM" eventid="1123" heatid="40040" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:02:47.40" entrycourse="SCM" eventid="1163" heatid="40121" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:01:20.37" entrycourse="SCM" eventid="1227" heatid="40203" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:30.94" entrycourse="SCM" eventid="1327" heatid="40383" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:00:36.84" entrycourse="SCM" eventid="1367" heatid="40449" lane="6">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Suchár" birthdate="2014-01-08" gender="M" nation="SVK" athleteid="38055">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.13" entrycourse="SCM" eventid="1133" heatid="40068" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:03:21.19" entrycourse="SCM" eventid="1153" heatid="40103" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:43.81" entrycourse="SCM" eventid="1173" heatid="40135" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:03:01.85" entrycourse="SCM" eventid="1197" heatid="40152" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:01:16.75" entrycourse="SCM" eventid="1237" heatid="40224" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:05:21.93" entrycourse="SCM" eventid="1257" heatid="40251" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:01:09.37" entrycourse="SCM" eventid="1277" heatid="40296" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:00:34.80" entrycourse="SCM" eventid="1297" heatid="40336" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:02:45.87" entrycourse="SCM" eventid="1317" heatid="40369" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:02:27.87" entrycourse="SCM" eventid="1357" heatid="40428" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:00:38.04" entrycourse="SCM" eventid="1377" heatid="40464" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:01:15.98" entrycourse="SCM" eventid="1397" heatid="40490" lane="3">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Barbora" lastname="Březnová" birthdate="2013-02-12" gender="F" nation="CZE" athleteid="38008">
              <ENTRIES>
                <ENTRY entrytime="00:02:56.38" entrycourse="SCM" eventid="1143" heatid="40098" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:37.07" entrycourse="SCM" eventid="1207" heatid="40172" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:11.15" entrycourse="SCM" eventid="1267" heatid="40271" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:01:18.10" entrycourse="SCM" eventid="1327" heatid="40390" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:42.06" entrycourse="SCM" eventid="1367" heatid="40441" lane="7">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alexej" lastname="Bátor" birthdate="2013-02-04" gender="M" nation="CZE" athleteid="37995">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.60" entrycourse="SCM" eventid="1133" heatid="40077" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:03:00.91" entrycourse="SCM" eventid="1153" heatid="40106" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:02:28.29" entrycourse="SCM" eventid="1173" heatid="40139" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:00:38.92" entrycourse="SCM" eventid="1217" heatid="40180" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:01:10.57" entrycourse="SCM" eventid="1237" heatid="40228" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:05:02.54" entrycourse="SCM" eventid="1257" heatid="40254" lane="2">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Klára" lastname="Pecová" birthdate="2012-11-16" gender="F" nation="CZE" athleteid="38047">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.19" entrycourse="SCM" eventid="1123" heatid="40038" lane="5">
                  <MEETINFO name="32. Int. Weihnachtsgala" city="Braunschweig" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:00:33.27" />
                </ENTRY>
                <ENTRY entrytime="00:03:20.46" entrycourse="SCM" eventid="1143" heatid="40092" lane="5">
                  <MEETINFO name="32. Int. Weihnachtsgala" city="Braunschweig" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:03:28.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.79" entrycourse="SCM" eventid="1207" heatid="40161" lane="4">
                  <MEETINFO name="32. Int. Weihnachtsgala" city="Braunschweig" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:00:46.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.94" entrycourse="SCM" eventid="1227" heatid="40199" lane="8">
                  <MEETINFO name="32. Int. Weihnachtsgala" city="Braunschweig" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:01:27.11" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.74" entrycourse="SCM" eventid="1267" heatid="40267" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:35.15" entrycourse="SCM" eventid="1327" heatid="40381" lane="8">
                  <MEETINFO name="32. Int. Weihnachtsgala" city="Braunschweig" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:01:39.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.93" entrycourse="LCM" eventid="1367" heatid="40443" lane="1">
                  <MEETINFO name="32. Int. Weihnachtsgala" city="Braunschweig" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:00:40.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marie" lastname="Štíbrová" birthdate="2014-07-27" gender="F" nation="CZE" athleteid="38098">
              <ENTRIES>
                <ENTRY entrytime="00:09:58.69" entrycourse="SCM" eventid="1083" heatid="40011" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:00:30.43" entrycourse="SCM" eventid="1123" heatid="40048" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:02:34.42" entrycourse="SCM" eventid="1163" heatid="40126" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:01:11.04" entrycourse="SCM" eventid="1227" heatid="40211" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:04:50.51" entrycourse="SCM" eventid="1247" heatid="40244" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:01:04.43" entrycourse="SCM" eventid="1267" heatid="40281" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:16.96" entrycourse="SCM" eventid="1347" heatid="40419" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:34.43" entrycourse="SCM" eventid="1367" heatid="40454" lane="5">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Štíbr" birthdate="2012-10-24" gender="M" nation="CZE" athleteid="38090">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.85" entrycourse="SCM" eventid="1133" heatid="40073" lane="5">
                </ENTRY>
                <ENTRY entrytime="00:02:55.38" entrycourse="SCM" eventid="1173" heatid="40132" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:01:21.64" entrycourse="SCM" eventid="1237" heatid="40221" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:05:09.43" entrycourse="SCM" eventid="1257" heatid="40253" lane="7">
                </ENTRY>
                <ENTRY entrytime="00:01:04.96" entrycourse="SCM" eventid="1277" heatid="40300" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:02:22.37" entrycourse="SCM" eventid="1357" heatid="40430" lane="6">
                </ENTRY>
                <ENTRY entrytime="00:00:38.65" entrycourse="LCM" eventid="1377" heatid="40464" lane="1">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Varga" birthdate="2014-05-15" gender="M" nation="CZE" athleteid="38068">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.12" entrycourse="SCM" eventid="1133" heatid="40068" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:03:00.97" entrycourse="SCM" eventid="1173" heatid="40131" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:48.74" entrycourse="SCM" eventid="1217" heatid="40174" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:05:46.54" entrycourse="SCM" eventid="1257" heatid="40248" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:14.39" entrycourse="SCM" eventid="1277" heatid="40293" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:40.17" entrycourse="SCM" eventid="1297" heatid="40332" lane="2">
                </ENTRY>
                <ENTRY entrytime="00:00:40.39" entrycourse="SCM" eventid="1377" heatid="40462" lane="4">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5637" nation="GER" region="03" clubid="35360" name="Zehlendorfer TSV von 1888 e.V.">
          <ATHLETES>
            <ATHLETE firstname="Freya Theresia Marie" lastname="Richter" birthdate="2015-01-01" gender="F" nation="GER" license="500100" athleteid="35369">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.15" eventid="1123" heatid="40027" lane="2">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:38.15" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.71" eventid="1227" heatid="40192" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:31.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.62" eventid="1267" heatid="40262" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:24.62" />
                </ENTRY>
                <ENTRY entrytime="00:03:30.00" eventid="1307" heatid="40348" lane="3">
                  <MEETINFO name="22. Seepferdchen-Cup" city="Potsdam" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:03:33.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.75" eventid="1367" heatid="40439" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:44.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Isabella Lilly" lastname="Gotzmann" birthdate="2015-01-01" gender="F" nation="GER" license="500097" athleteid="35361">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.80" eventid="1123" heatid="40027" lane="5">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:36.80" />
                </ENTRY>
                <ENTRY entrytime="00:03:25.00" eventid="1163" heatid="40112" lane="4" />
                <ENTRY entrytime="00:00:49.99" eventid="1207" heatid="40157" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:49.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.74" eventid="1227" heatid="40192" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:30.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.05" eventid="1267" heatid="40262" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:18.99" />
                </ENTRY>
                <ENTRY entrytime="00:03:30.00" eventid="1307" heatid="40348" lane="6">
                  <MEETINFO name="22. Seepferdchen-Cup" city="Potsdam" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:03:15.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.07" eventid="1367" heatid="40440" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:42.56" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5753" nation="GER" region="12" clubid="39084" name="Dresdner Delphine e.V.">
          <ATHLETES>
            <ATHLETE firstname="Jasna" lastname="Hänig" birthdate="2013-01-01" gender="F" nation="GER" license="445403" athleteid="39151">
              <ENTRIES>
                <ENTRY entrytime="00:05:59.99" eventid="1063" heatid="39995" lane="3">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-26" qualificationtime="00:06:23.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.82" eventid="1123" heatid="40041" lane="5">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:31.82" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.55" eventid="1163" heatid="40119" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:51.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.77" eventid="1187" heatid="40149" lane="1">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:02:50.77" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.51" eventid="1267" heatid="40276" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:01:08.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.74" eventid="1287" heatid="40324" lane="7">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:32.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.49" eventid="1387" heatid="40482" lane="3">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:14.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nils" lastname="Sonnabend" birthdate="2014-01-01" gender="M" nation="GER" license="454545" athleteid="39199">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.33" eventid="1133" heatid="40066" lane="8">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:31.58" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.41" eventid="1173" heatid="40131" lane="3">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:03:00.41" />
                </ENTRY>
                <ENTRY entrytime="00:03:20.00" eventid="1197" heatid="40151" lane="5" />
                <ENTRY entrytime="00:01:21.67" eventid="1237" heatid="40221" lane="1">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:21.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.88" eventid="1297" heatid="40336" lane="6">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:33.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:46.64" eventid="1317" heatid="40369" lane="7">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:02:46.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.99" eventid="1377" heatid="40465" lane="6">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:36.98" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ondrej" lastname="Bens" birthdate="2012-01-01" gender="M" nation="CZE" license="498809" athleteid="39087">
              <ENTRIES>
                <ENTRY entrytime="00:18:31.68" eventid="1113" heatid="40025" lane="2">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:19:30.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.00" eventid="1133" heatid="40072" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:00:30.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.65" eventid="1173" heatid="40133" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:51.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.00" eventid="1217" heatid="40180" lane="2" />
                <ENTRY entrytime="00:04:44.69" eventid="1257" heatid="40256" lane="3">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:05:00.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.33" eventid="1277" heatid="40301" lane="3">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:05.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.04" eventid="1317" heatid="40368" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:02:50.04" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.92" eventid="1357" heatid="40433" lane="1">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:02:22.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maximilian" lastname="Gennerich" birthdate="2011-01-01" gender="M" nation="GER" license="423096" athleteid="39135">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.72" eventid="1133" heatid="40080" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:26.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.00" eventid="1197" heatid="40154" lane="7" />
                <ENTRY entrytime="00:04:42.16" eventid="1257" heatid="40257" lane="7">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:04:42.16" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.82" eventid="1277" heatid="40307" lane="4">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:58.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.90" eventid="1297" heatid="40341" lane="4">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:28.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.60" eventid="1357" heatid="40435" lane="7">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-25" qualificationtime="00:02:10.60" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.45" eventid="1397" heatid="40494" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:02.96" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Milene" lastname="Müller" birthdate="2012-01-01" gender="F" nation="GER" license="437414" athleteid="39173">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.80" eventid="1123" heatid="40051" lane="1">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:00:29.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.53" eventid="1207" heatid="40171" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:37.05" />
                </ENTRY>
                <ENTRY entrytime="00:05:13.71" eventid="1247" heatid="40241" lane="2">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:05:13.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.12" eventid="1287" heatid="40322" lane="4">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:00:33.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.83" eventid="1327" heatid="40388" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:21.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.62" eventid="1387" heatid="40480" lane="5">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:17.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hannah" lastname="Böhmert" birthdate="2014-01-01" gender="F" nation="GER" license="447997" athleteid="39110">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.92" eventid="1123" heatid="40036" lane="8">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:32.05" />
                </ENTRY>
                <ENTRY entrytime="00:03:28.41" eventid="1143" heatid="40091" lane="2">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:03:28.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.91" eventid="1207" heatid="40163" lane="6">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:41.91" />
                </ENTRY>
                <ENTRY entrytime="00:05:44.82" eventid="1247" heatid="40236" lane="6">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:05:44.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.42" eventid="1267" heatid="40271" lane="1">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:11.42" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.76" eventid="1307" heatid="40355" lane="5">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:02:49.94" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.00" eventid="1347" heatid="40412" lane="1">
                  <MEETINFO name="Giraffenpokal" city="Chemnitz" course="LCM" approved="GER" date="2025-11-08" qualificationtime="00:02:34.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Kristof" lastname="Wagner" birthdate="2009-01-01" gender="M" nation="GER" license="395283" athleteid="39216">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.02" eventid="1133" heatid="40088" lane="1">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:25.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.04" eventid="1297" heatid="40346" lane="7">
                  <MEETINFO name="35. Herbstschwimmfest Zwickau" city="Zwickau" course="LCM" approved="GER" date="2025-11-15" qualificationtime="00:00:27.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Charlotte Katrin" lastname="Böhmert" birthdate="2013-01-01" gender="F" nation="GER" license="437495" athleteid="39096">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.28" eventid="1123" heatid="40034" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:32.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.75" eventid="1207" heatid="40160" lane="4">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:43.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.75" eventid="1227" heatid="40197" lane="4">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:24.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.78" eventid="1267" heatid="40269" lane="2">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:01:12.78" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.19" eventid="1307" heatid="40352" lane="6">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-27" qualificationtime="00:02:58.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.46" eventid="1367" heatid="40446" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:38.46" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Louis" lastname="Dramm" birthdate="2002-01-01" gender="M" nation="GER" license="282220" athleteid="39118">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.14" eventid="1133" heatid="40089" lane="2" />
                <ENTRY entrytime="00:00:50.20" eventid="1277" heatid="40311" lane="4">
                  <MEETINFO name="136. Deutsche Meisterschaften im Schwimmen" city="Berlin" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:00:50.20" />
                </ENTRY>
                <ENTRY entrytime="00:02:00.09" eventid="1317" heatid="40376" lane="4">
                  <MEETINFO name="136. Deutsche Meisterschaften im Schwimmen" city="Berlin" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:00.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.81" eventid="1397" heatid="40497" lane="4">
                  <MEETINFO name="136. Deutsche Meisterschaften im Schwimmen" city="Berlin" course="LCM" approved="GER" date="2025-05-01" qualificationtime="00:00:53.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marie-Sophie" lastname="Richter" birthdate="2014-01-01" gender="F" nation="GER" license="447792" athleteid="39180">
              <ENTRIES>
                <ENTRY entrytime="00:06:09.99" eventid="1063" heatid="39994" lane="6">
                  <MEETINFO name="Bezirksmeisterschaften Lange Strecke" city="Chemnitz" course="LCM" approved="GER" date="2025-01-26" qualificationtime="00:06:29.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.11" eventid="1123" heatid="40035" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:32.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:57.92" eventid="1163" heatid="40116" lane="4">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:02:57.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.63" eventid="1207" heatid="40165" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:39.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.35" eventid="1287" heatid="40320" lane="8">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:34.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.97" eventid="1327" heatid="40385" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:25.73" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.01" eventid="1347" heatid="40409" lane="3">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:40.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Luca" lastname="Egger" birthdate="2015-01-01" gender="M" nation="GER" license="463555" athleteid="39123">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.34" eventid="1133" heatid="40061" lane="3">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:36.00" />
                </ENTRY>
                <ENTRY entrytime="00:03:15.11" eventid="1173" heatid="40129" lane="3">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:03:15.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:49.68" eventid="1217" heatid="40174" lane="6">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:48.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.29" eventid="1237" heatid="40217" lane="6">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:29.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.40" eventid="1277" heatid="40291" lane="4">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:16.40" />
                </ENTRY>
                <ENTRY entrytime="00:03:02.96" eventid="1317" heatid="40365" lane="8">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:03:01.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.69" eventid="1377" heatid="40462" lane="1">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:40.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Vanessa" lastname="Illmann" birthdate="2002-01-01" gender="F" nation="GER" license="312872" athleteid="39224" />
            <ATHLETE firstname="Anna" lastname="Henze" birthdate="2013-01-01" gender="F" nation="GER" license="445341" athleteid="39159">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.31" eventid="1123" heatid="40053" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:28.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.66" eventid="1163" heatid="40123" lane="8">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:02:42.66" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.38" eventid="1227" heatid="40209" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:09.40" />
                </ENTRY>
                <ENTRY entrytime="00:05:08.19" eventid="1247" heatid="40242" lane="3">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:05:08.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.00" eventid="1267" heatid="40282" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:02.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.98" eventid="1367" heatid="40455" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:33.08" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.80" eventid="1387" heatid="40481" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:11.85" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Richard" lastname="Grohmann" birthdate="2001-01-01" gender="M" nation="GER" license="255122" athleteid="39223" />
            <ATHLETE firstname="Emil" lastname="Müller" birthdate="2009-01-01" gender="M" nation="GER" license="395288" athleteid="39167">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.18" eventid="1133" heatid="40085" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:25.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.70" eventid="1173" heatid="40141" lane="2">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:02:19.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.14" eventid="1277" heatid="40310" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:54.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.51" eventid="1317" heatid="40375" lane="2">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:02:21.51" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.80" eventid="1357" heatid="40437" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:57.46" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Matthäus" lastname="Haberkorn" birthdate="2012-01-01" gender="M" nation="GER" license="437400" athleteid="39143">
              <ENTRIES>
                <ENTRY entrytime="00:09:27.51" eventid="1093" heatid="40018" lane="2">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-12" qualificationtime="00:09:27.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.22" eventid="1133" heatid="40078" lane="4">
                  <MEETINFO name="29. Internationaler Plüschtierpokal" city="Dresden" course="LCM" approved="GER" date="2025-09-28" qualificationtime="00:00:28.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.04" eventid="1217" heatid="40184" lane="7">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:35.16" />
                </ENTRY>
                <ENTRY entrytime="00:04:41.07" eventid="1257" heatid="40257" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:04:32.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.12" eventid="1317" heatid="40372" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:25.20" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.25" eventid="1357" heatid="40433" lane="3">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:02:08.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.60" eventid="1397" heatid="40490" lane="1">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:09.34" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Niko" lastname="Srb" birthdate="2013-01-01" gender="M" nation="CZE" license="498813" athleteid="39207">
              <ENTRIES>
                <ENTRY entrytime="00:20:56.38" eventid="1113" heatid="40023" lane="5" />
                <ENTRY entrytime="00:00:34.40" eventid="1133" heatid="40064" lane="7">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:35.14" />
                </ENTRY>
                <ENTRY entrytime="00:03:19.53" eventid="1153" heatid="40103" lane="4">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-15" qualificationtime="00:03:31.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.37" eventid="1217" heatid="40178" lane="5">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:46.37" />
                </ENTRY>
                <ENTRY entrytime="00:05:23.33" eventid="1257" heatid="40251" lane="8">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:05:34.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.97" eventid="1277" heatid="40294" lane="8">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:15.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.96" eventid="1317" heatid="40365" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:03:09.94" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.47" eventid="1357" heatid="40425" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:42.02" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Flinn Jan" lastname="Böhmert" birthdate="2013-01-01" gender="M" nation="GER" license="437496" athleteid="39103">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.77" eventid="1133" heatid="40069" lane="5">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:31.77" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.97" eventid="1173" heatid="40134" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:02:49.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.39" eventid="1237" heatid="40223" lane="6">
                  <MEETINFO name="33. Internationale Geraer Stadtmeisterschaften" city="Gera" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:18.39" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.36" eventid="1277" heatid="40295" lane="4">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:10.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.23" eventid="1297" heatid="40335" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:35.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.41" eventid="1357" heatid="40424" lane="5">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:02:39.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Liesbeth" lastname="Sauer" birthdate="2012-01-01" gender="F" nation="GER" license="444965" athleteid="39188">
              <ENTRIES>
                <ENTRY entrytime="00:02:58.38" eventid="1143" heatid="40098" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:58.38" />
                </ENTRY>
                <ENTRY entrytime="00:05:18.11" eventid="1247" heatid="40240" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:05:18.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.11" eventid="1287" heatid="40327" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:30.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.46" eventid="1327" heatid="40389" lane="5">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:01:20.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.13" eventid="1367" heatid="40453" lane="2">
                  <MEETINFO name="14. Internationales Sprintmeeting des OSSV Kamenz" city="Kamenz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.85" eventid="1387" heatid="40483" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:10.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alina" lastname="Zubovska" birthdate="2009-01-01" gender="F" nation="UKR" license="454879" athleteid="39219">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.39" eventid="1287" heatid="40329" lane="7">
                  <MEETINFO name="Kinder- und Jugendspiele der Stadt Dresden" city="Dresden" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:00:29.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.94" eventid="1367" heatid="40459" lane="1">
                  <MEETINFO name="10. Dresdner Elbepokal" city="Dresden" course="LCM" approved="GER" date="2025-09-14" qualificationtime="00:00:31.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lennard" lastname="Barthel" birthdate="2013-01-01" gender="M" nation="GER" license="437409" athleteid="39085">
              <ENTRIES>
                <ENTRY entrytime="00:20:05.31" eventid="1113" heatid="40024" lane="2">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:23:05.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Engel" birthdate="2001-01-01" gender="M" nation="GER" license="256573" athleteid="39131">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.29" eventid="1297" heatid="40347" lane="3">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:00:25.27" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marlin" lastname="Garsuch" birthdate="2004-01-01" gender="F" nation="GER" license="315358" athleteid="39133">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.40" eventid="1123" heatid="40056" lane="8">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-31" qualificationtime="00:00:28.40" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Schaarschmidt" birthdate="2003-01-01" gender="F" nation="GER" license="297766" athleteid="39195">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.59" eventid="1123" heatid="40052" lane="7">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-31" qualificationtime="00:00:29.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.00" eventid="1267" heatid="40273" lane="1" />
                <ENTRY entrytime="00:02:54.74" eventid="1307" heatid="40354" lane="8">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-07" qualificationtime="00:02:54.74" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Amadeus" lastname="Bräuning" birthdate="1998-01-01" gender="M" nation="GER" license="173989" athleteid="39222" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.00" eventid="1185" heatid="40146" lane="6">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" date="2025-06-15" qualificationtime="00:01:53.48" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.85" eventid="1185" heatid="40146" lane="2">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" date="2025-06-15" qualificationtime="00:01:53.48" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.00" eventid="1183" heatid="40144" lane="6">
                  <MEETINFO name="47. Schwimmzonen- und Mastersmeeting" city="Enns" date="2025-06-15" qualificationtime="00:02:08.63" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="3386" nation="GER" region="12" clubid="38846" name="SV Dresden-Nord">
          <ATHLETES>
            <ATHLETE firstname="Cara" lastname="Noeske" birthdate="2011-01-01" gender="F" nation="GER" license="436299" athleteid="38849">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.82" eventid="1123" heatid="40033" lane="1">
                  <MEETINFO name="6. Frühjahrswettkampf" city="Dresden" course="SCM" approved="GER" date="2025-03-23" qualificationtime="00:00:33.82" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Böhme" birthdate="2010-01-01" gender="M" nation="GER" license="511851" athleteid="38847">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.42" eventid="1133" heatid="40072" lane="1">
                  <MEETINFO name="6. Herbstwettkampf der SG EDM" city="Dresden" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:00:30.42" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Martin" lastname="Schmidt" birthdate="2008-01-01" gender="M" nation="GER" license="379866" athleteid="38860">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.23" eventid="1277" heatid="40303" lane="1">
                  <MEETINFO name="26. Internationaler WTC-Pokal" city="Dresden" course="LCM" approved="GER" date="2025-12-06" qualificationtime="00:01:02.23" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Max" lastname="Olbrich" birthdate="2014-01-01" gender="M" nation="GER" license="474578" athleteid="38851">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.96" eventid="1133" heatid="40062" lane="8">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:35.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.12" eventid="1217" heatid="40177" lane="3">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:44.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.77" eventid="1277" heatid="40288" lane="7">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:24.77" />
                </ENTRY>
                <ENTRY entrytime="00:01:39.81" eventid="1337" heatid="40392" lane="4">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:39.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Amelie" lastname="Podworny" birthdate="2010-01-01" gender="F" nation="GER" license="410084" athleteid="38856">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.66" eventid="1123" heatid="40030" lane="4">
                  <MEETINFO name="6. Herbstwettkampf der SG EDM" city="Dresden" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:00:34.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Malte" lastname="Progscha" birthdate="2012-01-01" gender="M" nation="GER" license="449960" athleteid="38858">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.97" eventid="1133" heatid="40063" lane="1">
                  <MEETINFO name="6. Herbstwettkampf der SG EDM" city="Dresden" course="LCM" approved="GER" date="2025-11-09" qualificationtime="00:00:34.97" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3261" nation="GER" region="16" clubid="37124" name="SV Nordhausen 90 e.V.">
          <ATHLETES>
            <ATHLETE firstname="Frida" lastname="Flagmeyer" birthdate="2014-01-01" gender="F" nation="GER" license="448053" athleteid="38916">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.18" eventid="1123" heatid="40039" lane="8">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:32.18" />
                </ENTRY>
                <ENTRY entrytime="00:03:17.39" eventid="1143" heatid="40093" lane="7">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:03:17.39" />
                </ENTRY>
                <ENTRY entrytime="00:03:00.06" eventid="1187" heatid="40148" lane="7">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:03:00.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.35" eventid="1287" heatid="40320" lane="1">
                  <MEETINFO name="31. off Landesmeisterschaften mit JG-u Kindermeist" city="Magdeburg" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:34.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.90" eventid="1327" heatid="40382" lane="7">
                  <MEETINFO name="Überprüfungswettkampf" city="Halle (Saale)" course="LCM" approved="GER" date="2025-02-07" qualificationtime="00:01:31.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Tom" lastname="Falke" birthdate="2010-01-01" gender="M" nation="GER" license="397841" athleteid="38910">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.48" eventid="1133" heatid="40078" lane="8">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:28.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.39" eventid="1217" heatid="40183" lane="3">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:35.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.44" eventid="1297" heatid="40336" lane="4">
                  <MEETINFO name="Dresdner Tage der Talente" city="Dresden" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:00:33.44" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.44" eventid="1317" heatid="40370" lane="1">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:02:44.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.22" eventid="1377" heatid="40468" lane="6">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:34.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Karl-Justus" lastname="Höpfner" birthdate="2013-01-01" gender="M" nation="GER" license="442342" athleteid="38922">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.99" eventid="1277" heatid="40289" lane="4">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:15.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.95" eventid="1297" heatid="40332" lane="4">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:37.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.35" eventid="1337" heatid="40393" lane="4">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:30.69" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.16" eventid="1397" heatid="40487" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:01:31.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="37136" firstname="Paul-Emil" gender="M" grade="WKR" lastname="Höpfner" nation="GER" />
            <OFFICIAL officialid="38927" firstname="Paul-Emil" gender="M" grade="WKR" lastname="Höpfner" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="2502" nation="GER" region="18" clubid="35169" name="SV Cannstatt">
          <ATHLETES>
            <ATHLETE firstname="Matilda" lastname="Biedermann" birthdate="2013-01-01" gender="F" nation="GER" license="457104" athleteid="37632">
              <ENTRIES>
                <ENTRY entrytime="00:06:05.48" eventid="1063" heatid="39995" lane="1">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:06:05.48" />
                </ENTRY>
                <ENTRY entrytime="00:03:12.33" eventid="1143" heatid="40094" lane="7">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:03:02.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.27" eventid="1207" heatid="40164" lane="5">
                  <MEETINFO name="BaWü-Jahrgangsmeisterschaften (jüngere Jahrgänge)" city="Heidelberg" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:00:41.27" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.66" eventid="1227" heatid="40195" lane="6">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:23.98" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.43" eventid="1307" heatid="40351" lane="2">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:52.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.97" eventid="1327" heatid="40382" lane="8">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:28.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.05" eventid="1347" heatid="40407" lane="7">
                  <MEETINFO name="SUN-RISE Meeting" city="Neckarsulm" course="LCM" approved="GER" date="2025-02-02" qualificationtime="00:02:50.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Josef" lastname="Mittermeier" birthdate="2012-01-01" gender="M" nation="GER" license="445919" athleteid="37727">
              <ENTRIES>
                <ENTRY entrytime="00:10:29.00" eventid="1093" heatid="40016" lane="8">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-09" qualificationtime="00:10:47.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.98" eventid="1133" heatid="40071" lane="1">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:30.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.47" eventid="1173" heatid="40134" lane="4">
                  <MEETINFO name="8. Backnanger Schwimmfest" city="Backnang" course="SCM" approved="GER" date="2025-05-03" qualificationtime="00:02:44.39" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.03" eventid="1237" heatid="40221" lane="5">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:17.78" />
                </ENTRY>
                <ENTRY entrytime="00:05:08.82" eventid="1257" heatid="40253" lane="2">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:05:05.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.21" eventid="1277" heatid="40298" lane="7">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:06.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.59" eventid="1317" heatid="40367" lane="7">
                  <MEETINFO name="SV Cannstatt Young Challenge" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-10-05" qualificationtime="00:02:47.35" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.45" eventid="1357" heatid="40429" lane="8">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:22.56" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lia" lastname="Laschinsky" birthdate="2008-01-01" gender="F" nation="GER" license="365049" athleteid="37795">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.59" eventid="1123" heatid="40052" lane="2">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:00:29.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.36" eventid="1163" heatid="40125" lane="1">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-10" qualificationtime="00:02:39.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.36" eventid="1227" heatid="40210" lane="4">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:01:10.08" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.14" eventid="1267" heatid="40280" lane="4">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:01:05.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.36" eventid="1287" heatid="40327" lane="2">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:00:31.36" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.71" eventid="1347" heatid="40416" lane="2">
                  <MEETINFO name="Württembergische Meisterschaften" city="Böblingen" course="LCM" approved="GER" date="2025-07-19" qualificationtime="00:02:25.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.65" eventid="1367" heatid="40458" lane="8">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-23" qualificationtime="00:00:32.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Franziska" lastname="Maier" birthdate="2012-01-01" gender="F" nation="GER" license="439715" athleteid="37709">
              <ENTRIES>
                <ENTRY entrytime="00:10:28.00" eventid="1083" heatid="40009" lane="3">
                  <MEETINFO name="Ba-Wü Meisterschaften Lange Strecke incl. Masters" city="Karlsruhe" course="LCM" approved="GER" date="2025-02-08" qualificationtime="00:11:18.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.08" eventid="1123" heatid="40045" lane="2">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:30.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.83" eventid="1163" heatid="40120" lane="3">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:44.21" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.55" eventid="1227" heatid="40204" lane="7">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:15.42" />
                </ENTRY>
                <ENTRY entrytime="00:05:20.83" eventid="1247" heatid="40239" lane="1">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:05:11.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.47" eventid="1267" heatid="40276" lane="5">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:07.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.30" eventid="1287" heatid="40317" lane="3">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:33.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.92" eventid="1347" heatid="40414" lane="8">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:27.33" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Wetzlberger" birthdate="2013-01-01" gender="F" nation="GER" license="467534" athleteid="37754">
              <ENTRIES>
                <ENTRY entrytime="00:06:09.00" eventid="1063" heatid="39994" lane="5">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-09" qualificationtime="00:06:22.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.92" eventid="1123" heatid="40032" lane="3">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:32.74" />
                </ENTRY>
                <ENTRY entrytime="00:03:06.45" eventid="1163" heatid="40114" lane="4">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:51.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.68" eventid="1207" heatid="40162" lane="7">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:42.68" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.61" eventid="1227" heatid="40196" lane="1">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:20.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.41" eventid="1267" heatid="40267" lane="6">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:13.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.12" eventid="1307" heatid="40352" lane="1">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:54.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.84" eventid="1347" heatid="40409" lane="8">
                  <MEETINFO name="BaWü &amp; Süddt Meisterschaften SMK" city="Stuttgart" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:41.84" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Zahn" birthdate="2013-01-01" gender="M" nation="GER" license="476703" athleteid="37763">
              <ENTRIES>
                <ENTRY entrytime="00:10:35.00" eventid="1093" heatid="40015" lane="2">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-09" qualificationtime="00:11:15.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.39" eventid="1133" heatid="40072" lane="7">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:29.85" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.79" eventid="1173" heatid="40134" lane="6">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:44.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.54" eventid="1217" heatid="40177" lane="4">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:43.54" />
                </ENTRY>
                <ENTRY entrytime="00:05:25.64" eventid="1257" heatid="40250" lane="3">
                  <MEETINFO name="BaWü-Jahrgangsmeisterschaften (jüngere Jahrgänge)" city="Heidelberg" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:05:25.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.90" eventid="1277" heatid="40297" lane="6">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:01:07.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:57.69" eventid="1317" heatid="40366" lane="1">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:44.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.29" eventid="1357" heatid="40427" lane="2">
                  <MEETINFO name="BaWü &amp; Süddt Meisterschaften SMK" city="Stuttgart" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:32.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Tim" lastname="Sauer" birthdate="2008-01-01" gender="M" nation="GER" license="403613" athleteid="37803">
              <ENTRIES>
                <ENTRY entrytime="00:09:33.47" eventid="1093" heatid="40018" lane="8">
                  <MEETINFO name="58. ISTKa" city="Karlsruhe" course="LCM" approved="GER" date="2025-12-05" qualificationtime="00:09:09.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.45" eventid="1133" heatid="40084" lane="5">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-29" qualificationtime="00:00:26.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.62" eventid="1197" heatid="40154" lane="4">
                  <MEETINFO name="Ba-Wü Meisterschaften Lange Strecke incl. Masters" city="Karlsruhe" course="LCM" approved="GER" date="2025-02-08" qualificationtime="00:02:26.62" />
                </ENTRY>
                <ENTRY entrytime="00:04:23.88" eventid="1257" heatid="40259" lane="7">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:04:23.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.45" eventid="1277" heatid="40310" lane="2">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:54.99" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.76" eventid="1317" heatid="40375" lane="7">
                  <MEETINFO name="SV Cannstatt Young Challenge" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-10-05" qualificationtime="00:02:19.96" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.31" eventid="1357" heatid="40438" lane="2">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:00.02" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Regina" lastname="Meintzinger" birthdate="2013-01-01" gender="F" nation="GER" license="452141" athleteid="37718">
              <ENTRIES>
                <ENTRY entrytime="00:11:27.08" eventid="1083" heatid="40005" lane="5">
                  <MEETINFO name="20. Schwaben-Cup" city="Stuttgart" course="LCM" approved="GER" date="2025-04-04" qualificationtime="00:11:27.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.04" eventid="1123" heatid="40035" lane="6">
                  <MEETINFO name="Swim Race Days Dortmund" city="Dortmund" course="LCM" approved="GER" date="2025-03-01" qualificationtime="00:00:33.04" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.15" eventid="1163" heatid="40118" lane="3">
                  <MEETINFO name="BaWü-Jahrgangsmeisterschaften (jüngere Jahrgänge)" city="Heidelberg" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:02:53.15" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.04" eventid="1227" heatid="40198" lane="4">
                  <MEETINFO name="BaWü-Jahrgangsmeisterschaften (jüngere Jahrgänge)" city="Heidelberg" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:20.73" />
                </ENTRY>
                <ENTRY entrytime="00:05:31.13" eventid="1247" heatid="40237" lane="5">
                  <MEETINFO name="Ba-Wü Meisterschaften Lange Strecke incl. Masters" city="Karlsruhe" course="LCM" approved="GER" date="2025-02-09" qualificationtime="00:05:31.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.20" eventid="1267" heatid="40270" lane="2">
                  <MEETINFO name="Swim Race Days Dortmund" city="Dortmund" course="LCM" approved="GER" date="2025-03-02" qualificationtime="00:01:12.20" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.18" eventid="1307" heatid="40354" lane="7">
                  <MEETINFO name="BaWü &amp; Süddt Meisterschaften SMK" city="Stuttgart" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:54.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.17" eventid="1347" heatid="40410" lane="7">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:35.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lui Luke" lastname="Aderhold" birthdate="2013-01-01" gender="M" nation="GER" license="454320" athleteid="37623">
              <ENTRIES>
                <ENTRY entrytime="00:10:44.00" eventid="1093" heatid="40014" lane="5">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-09" qualificationtime="00:11:18.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.57" eventid="1133" heatid="40067" lane="4">
                  <MEETINFO name="SV Cannstatt Young Challenge" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-10-05" qualificationtime="00:00:31.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.23" eventid="1173" heatid="40133" lane="8">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:46.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.98" eventid="1237" heatid="40222" lane="6">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:17.33" />
                </ENTRY>
                <ENTRY entrytime="00:05:27.99" eventid="1257" heatid="40250" lane="8">
                  <MEETINFO name="BaWü &amp; Süddt Meisterschaften SMK" city="Stuttgart" course="LCM" approved="GER" date="2025-05-02" qualificationtime="00:05:27.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.08" eventid="1277" heatid="40296" lane="1">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-28" qualificationtime="00:01:10.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:58.06" eventid="1317" heatid="40366" lane="8">
                  <MEETINFO name="BaWü &amp; Süddt Meisterschaften SMK" city="Stuttgart" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:02:58.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.79" eventid="1357" heatid="40425" lane="7">
                  <MEETINFO name="8. Backnanger Schwimmfest" city="Backnang" course="SCM" approved="GER" date="2025-05-03" qualificationtime="00:02:37.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Rieke" lastname="Blümel" birthdate="2012-01-01" gender="F" nation="GER" license="437297" athleteid="37640">
              <ENTRIES>
                <ENTRY entrytime="00:10:40.96" eventid="1083" heatid="40009" lane="7">
                  <MEETINFO name="Challenge Jacky Ernewein" city="Strasbourg" course="LCM" approved="GER" date="2025-01-24" qualificationtime="00:10:40.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.90" eventid="1123" heatid="40050" lane="5">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:28.82" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.11" eventid="1163" heatid="40125" lane="6">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:31.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.05" eventid="1187" heatid="40150" lane="1">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:36.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.71" eventid="1227" heatid="40210" lane="2">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:08.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.90" eventid="1267" heatid="40282" lane="4">
                  <MEETINFO name="DMSJ Bundesfinale" city="Wuppertal" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:00.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.10" eventid="1307" heatid="40359" lane="5">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:34.29" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.32" eventid="1347" heatid="40417" lane="2">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-29" qualificationtime="00:02:23.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Aylan" lastname="Isougri" birthdate="2012-01-01" gender="M" nation="GER" license="431523" athleteid="37674">
              <ENTRIES>
                <ENTRY entrytime="00:10:30.00" eventid="1093" heatid="40015" lane="5" />
                <ENTRY entrytime="00:00:32.62" eventid="1133" heatid="40067" lane="3">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:31.57" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.38" eventid="1173" heatid="40132" lane="8">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:49.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.40" eventid="1237" heatid="40220" lane="2">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:22.18" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.65" eventid="1277" heatid="40294" lane="4">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:09.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.42" eventid="1337" heatid="40394" lane="6">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:29.80" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.43" eventid="1357" heatid="40426" lane="2">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:02:35.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Parsa" lastname="Ezadi" birthdate="2010-01-01" gender="M" nation="GER" license="482097" athleteid="37772">
              <ENTRIES>
                <ENTRY entrytime="00:10:21.31" eventid="1093" heatid="40016" lane="6" />
                <ENTRY entrytime="00:00:28.42" eventid="1133" heatid="40078" lane="1">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-29" qualificationtime="00:00:28.42" />
                </ENTRY>
                <ENTRY entrytime="00:04:56.56" eventid="1257" heatid="40255" lane="1">
                  <MEETINFO name="International Sindelfingen Swimming Championship" city="Sindelfingen" course="LCM" approved="GER" date="2025-03-22" qualificationtime="00:04:56.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.23" eventid="1277" heatid="40303" lane="8">
                  <MEETINFO name="SV Cannstatt Young Challenge" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-10-05" qualificationtime="00:01:01.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.06" eventid="1297" heatid="40337" lane="7">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-28" qualificationtime="00:00:33.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.63" eventid="1317" heatid="40371" lane="1">
                  <MEETINFO name="SV Cannstatt Young Challenge" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-10-05" qualificationtime="00:02:34.93" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.70" eventid="1357" heatid="40431" lane="2">
                  <MEETINFO name="International Sindelfingen Swimming Championship" city="Sindelfingen" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:02:18.70" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Franziska" lastname="Grimm" birthdate="2013-01-01" gender="F" nation="GER" license="447098" athleteid="37658">
              <ENTRIES>
                <ENTRY entrytime="00:11:14.00" eventid="1083" heatid="40006" lane="2">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-09" qualificationtime="00:11:44.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.64" eventid="1123" heatid="40029" lane="1">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:34.99" />
                </ENTRY>
                <ENTRY entrytime="00:03:07.82" eventid="1143" heatid="40095" lane="2">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:03:03.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.31" eventid="1207" heatid="40164" lane="3">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:40.46" />
                </ENTRY>
                <ENTRY entrytime="00:03:02.61" eventid="1307" heatid="40351" lane="3">
                  <MEETINFO name="Württembergische Meisterschaften" city="Böblingen" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:03:02.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.65" eventid="1327" heatid="40384" lane="4">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:26.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.15" eventid="1347" heatid="40408" lane="8">
                  <MEETINFO name="20. Schwaben-Cup" city="Stuttgart" course="LCM" approved="GER" date="2025-04-06" qualificationtime="00:02:45.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Eleni" lastname="Kementzetzidou" birthdate="2013-01-01" gender="F" nation="GER" license="452342" athleteid="37691">
              <ENTRIES>
                <ENTRY entrytime="00:06:00.92" eventid="1063" heatid="39995" lane="2">
                  <MEETINFO name="SV Cannstatt Überprüfungswettkampf" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:05:46.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.55" eventid="1123" heatid="40034" lane="8" />
                <ENTRY entrytime="00:02:43.86" eventid="1163" heatid="40122" lane="6">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:41.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.77" eventid="1207" heatid="40171" lane="1">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:37.05" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.42" eventid="1227" heatid="40208" lane="1">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:13.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.65" eventid="1287" heatid="40321" lane="3">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:32.24" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.23" eventid="1307" heatid="40357" lane="1">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:40.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.79" eventid="1347" heatid="40412" lane="2">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:02:33.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Sommerlatte" birthdate="2012-01-01" gender="M" nation="GER" license="445864" athleteid="37736">
              <ENTRIES>
                <ENTRY entrytime="00:05:18.67" eventid="1073" heatid="40001" lane="1">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:05:03.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.35" eventid="1133" heatid="40075" lane="6">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:28.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.01" eventid="1153" heatid="40110" lane="1">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:35.42" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.65" eventid="1197" heatid="40154" lane="8">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:31.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.83" eventid="1217" heatid="40184" lane="4">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:00:35.83" />
                </ENTRY>
                <ENTRY entrytime="00:04:45.48" eventid="1257" heatid="40256" lane="7">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:04:35.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.92" eventid="1317" heatid="40372" lane="6">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:02:25.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.87" eventid="1337" heatid="40401" lane="8">
                  <MEETINFO name="DMSJ Württemberg-Finale" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:11.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.16" eventid="1357" heatid="40432" lane="8">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:13.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lina" lastname="Hellenthal" birthdate="2011-01-01" gender="F" nation="GER" license="432636" athleteid="37780">
              <ENTRIES>
                <ENTRY entrytime="00:10:46.98" eventid="1083" heatid="40008" lane="3">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-09" qualificationtime="00:10:46.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.82" eventid="1163" heatid="40117" lane="3">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-10" qualificationtime="00:02:55.82" />
                </ENTRY>
                <ENTRY entrytime="00:05:13.26" eventid="1247" heatid="40241" lane="3">
                  <MEETINFO name="20. Internationaler Bären – Cup" city="Waldenbuch" course="SCM" approved="GER" date="2025-10-04" qualificationtime="00:05:12.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.79" eventid="1267" heatid="40271" lane="8">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-28" qualificationtime="00:01:11.79" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.12" eventid="1307" heatid="40354" lane="4">
                  <MEETINFO name="SV Cannstatt Young Challenge" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-10-05" qualificationtime="00:02:51.99" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.83" eventid="1347" heatid="40412" lane="7">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-29" qualificationtime="00:02:34.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Johannes" lastname="Weeger" birthdate="2010-01-01" gender="M" nation="GER" license="411846" athleteid="37811">
              <ENTRIES>
                <ENTRY entrytime="00:05:05.59" eventid="1073" heatid="40001" lane="2">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-17" qualificationtime="00:04:51.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.05" eventid="1133" heatid="40083" lane="8">
                  <MEETINFO name="41. AchalmCup" city="Reutlingen" course="LCM" approved="GER" date="2025-06-29" qualificationtime="00:00:27.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.20" eventid="1153" heatid="40109" lane="1">
                  <MEETINFO name="Württembergische Meisterschaften" city="Böblingen" course="LCM" approved="GER" date="2025-07-20" qualificationtime="00:02:47.20" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.97" eventid="1197" heatid="40155" lane="2">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:02:21.97" />
                </ENTRY>
                <ENTRY entrytime="00:04:38.41" eventid="1257" heatid="40258" lane="7">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:04:27.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.70" eventid="1277" heatid="40308" lane="7">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:57.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.37" eventid="1317" heatid="40374" lane="8">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:19.26" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.54" eventid="1357" heatid="40434" lane="4">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:02:11.54" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Neo" lastname="Engelmann" birthdate="2013-01-01" gender="M" nation="GER" license="446819" athleteid="37649">
              <ENTRIES>
                <ENTRY entrytime="00:10:44.00" eventid="1093" heatid="40014" lane="3">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-09" qualificationtime="00:11:07.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.16" eventid="1133" heatid="40066" lane="6">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:32.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.99" eventid="1173" heatid="40134" lane="7">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:41.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.17" eventid="1237" heatid="40221" lane="6">
                  <MEETINFO name="DMSJ Württemberg-Finale" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-11-23" qualificationtime="00:01:14.68" />
                </ENTRY>
                <ENTRY entrytime="00:05:22.61" eventid="1257" heatid="40251" lane="1">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:05:15.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.03" eventid="1277" heatid="40294" lane="6">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:11.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.61" eventid="1317" heatid="40366" lane="3">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:47.80" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.83" eventid="1357" heatid="40426" lane="5">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:29.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilia Sophia" lastname="Zeh" birthdate="2007-01-01" gender="F" nation="GER" license="402397" athleteid="37820">
              <ENTRIES>
                <ENTRY entrytime="00:05:10.98" eventid="1063" heatid="39997" lane="6">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-17" qualificationtime="00:05:01.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.56" eventid="1143" heatid="40099" lane="2">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:02:40.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.47" eventid="1207" heatid="40173" lane="8">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-10" qualificationtime="00:00:36.16" />
                </ENTRY>
                <ENTRY entrytime="00:04:38.28" eventid="1247" heatid="40245" lane="2">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:04:32.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.05" eventid="1287" heatid="40328" lane="2">
                  <MEETINFO name="International Sindelfingen Swimming Championship" city="Sindelfingen" course="LCM" approved="GER" date="2025-03-22" qualificationtime="00:00:31.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.21" eventid="1327" heatid="40390" lane="3">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:14.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Yassir" lastname="Lahrach" birthdate="2013-01-01" gender="M" nation="GER" license="443497" athleteid="37700">
              <ENTRIES>
                <ENTRY entrytime="00:06:01.03" eventid="1073" heatid="39999" lane="7">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-17" qualificationtime="00:05:29.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.24" eventid="1133" heatid="40072" lane="2">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:29.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.18" eventid="1173" heatid="40136" lane="8">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:35.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.58" eventid="1237" heatid="40223" lane="4">
                  <MEETINFO name="DMSJ Württemberg-Finale" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:12.81" />
                </ENTRY>
                <ENTRY entrytime="00:05:05.14" eventid="1257" heatid="40254" lane="8">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:04:57.39" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.66" eventid="1277" heatid="40299" lane="1">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:01:04.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.31" eventid="1317" heatid="40370" lane="5">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:34.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.75" eventid="1357" heatid="40430" lane="1">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:02:19.56" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ayman" lastname="Isougri" birthdate="2012-01-01" gender="M" nation="GER" license="431525" athleteid="37682">
              <ENTRIES>
                <ENTRY entrytime="00:10:30.00" eventid="1093" heatid="40015" lane="3" />
                <ENTRY entrytime="00:00:33.03" eventid="1133" heatid="40067" lane="8">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:32.64" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.66" eventid="1173" heatid="40132" lane="3">
                  <MEETINFO name="15. Internationaler Sendercup" city="Mühlacker" course="LCM" approved="GER" date="2025-06-01" qualificationtime="00:02:56.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.26" eventid="1217" heatid="40178" lane="4">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:42.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.45" eventid="1237" heatid="40220" lane="7">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:19.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.01" eventid="1277" heatid="40294" lane="3">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:11.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.37" eventid="1337" heatid="40395" lane="1">
                  <MEETINFO name="46. HEDINT" city="Heddesheim" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:01:32.37" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.50" eventid="1357" heatid="40425" lane="5">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:02:36.50" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Pia" lastname="Ketterer" birthdate="2009-01-01" gender="F" nation="GER" license="399365" athleteid="37787">
              <ENTRIES>
                <ENTRY entrytime="00:05:43.08" eventid="1063" heatid="39996" lane="6" />
                <ENTRY entrytime="00:00:29.69" eventid="1123" heatid="40051" lane="6">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-10" qualificationtime="00:00:30.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.17" eventid="1227" heatid="40206" lane="4">
                  <MEETINFO name="SV Cannstatt Young Challenge" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-10-05" qualificationtime="00:01:15.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.05" eventid="1287" heatid="40328" lane="7">
                  <MEETINFO name="73. Süddeutsche Meisterschaften offen u. Jahrgang" city="Stuttgart" course="LCM" approved="GER" date="2025-05-23" qualificationtime="00:00:31.17" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.25" eventid="1307" heatid="40358" lane="5">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:36.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.75" eventid="1347" heatid="40416" lane="7">
                  <MEETINFO name="Challenge Jacky Ernewein" city="Strasbourg" course="LCM" approved="GER" date="2025-01-25" qualificationtime="00:02:40.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.02" eventid="1367" heatid="40453" lane="5">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:00:35.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Moritz Peter" lastname="Grimm" birthdate="2012-01-01" gender="M" nation="GER" license="438235" athleteid="37666">
              <ENTRIES>
                <ENTRY entrytime="00:10:28.79" eventid="1093" heatid="40016" lane="1">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-09" qualificationtime="00:10:28.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.39" eventid="1133" heatid="40065" lane="4">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:33.06" />
                </ENTRY>
                <ENTRY entrytime="00:03:12.87" eventid="1153" heatid="40104" lane="5">
                  <MEETINFO name="International Sindelfingen Swimming Championship" city="Sindelfingen" course="LCM" approved="GER" date="2025-03-23" qualificationtime="00:03:12.87" />
                </ENTRY>
                <ENTRY entrytime="00:05:07.52" eventid="1257" heatid="40253" lane="3">
                  <MEETINFO name="Baden-Württembergische Kurzbahn-Meisterschaften" city="Neckarsulm" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:05:04.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.54" eventid="1317" heatid="40367" lane="5">
                  <MEETINFO name="8. Backnanger Schwimmfest" city="Backnang" course="SCM" approved="GER" date="2025-05-03" qualificationtime="00:02:46.66" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.37" eventid="1337" heatid="40395" lane="6">
                  <MEETINFO name="4. Internationales Feuerbacher Kurzbahnmeeting" city="Stuttgart" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:25.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.57" eventid="1357" heatid="40428" lane="2">
                  <MEETINFO name="49. International Dr. Otto-Fahr Swim-Meeting" city="Stuttgart" course="LCM" approved="GER" date="2025-05-11" qualificationtime="00:02:28.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="40501" name="Ustecka akademie plaveckych sportu" shortname="UAPS">
          <ATHLETES>
            <ATHLETE firstname="Janecek" lastname="Vojtech" birthdate="2001-01-01" gender="M" nation="CZE" athleteid="40502">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.52" eventid="1217" heatid="40190" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4743" nation="GER" region="04" clubid="36905" name="Neptun 08 Finsterwalde e.V.">
          <ATHLETES>
            <ATHLETE firstname="Fiona" lastname="Fröschke" birthdate="2010-01-01" gender="F" nation="GER" license="411635" athleteid="36914">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.02" eventid="1123" heatid="40046" lane="1">
                  <MEETINFO name="Schwimmfest zum Jahrestag der Schwimmhalle" city="Forst" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:30.85" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.41" eventid="1143" heatid="40098" lane="3">
                  <MEETINFO name="14. Sängerpokal" city="Finsterwalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:53.41" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.80" eventid="1163" heatid="40123" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:40.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.93" eventid="1207" heatid="40172" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:36.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.69" eventid="1227" heatid="40208" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:14.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.46" eventid="1287" heatid="40325" lane="7">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:00:32.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.85" eventid="1307" heatid="40358" lane="4">
                  <MEETINFO name="14. Sängerpokal" city="Finsterwalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:38.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.04" eventid="1327" heatid="40389" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:20.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Dean" lastname="Schöne" birthdate="2013-01-01" gender="M" nation="GER" license="446291" athleteid="36942">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.49" eventid="1133" heatid="40070" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:31.49" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.33" eventid="1153" heatid="40106" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:03:03.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.35" eventid="1217" heatid="40181" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:38.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.57" eventid="1237" heatid="40217" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:28.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.86" eventid="1277" heatid="40295" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:10.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.23" eventid="1297" heatid="40335" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:35.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.40" eventid="1317" heatid="40368" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:50.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.16" eventid="1337" heatid="40396" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:27.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lore" lastname="Kittler" birthdate="2015-01-01" gender="F" nation="GER" license="467147" athleteid="36932">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.66" eventid="1123" heatid="40026" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:39.66" />
                </ENTRY>
                <ENTRY entrytime="00:03:29.95" eventid="1163" heatid="40112" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:03:29.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.75" eventid="1227" heatid="40192" lane="2">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:37.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Georg" lastname="Gärtner" birthdate="2013-01-01" gender="M" nation="GER" license="446154" athleteid="36923">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.15" eventid="1133" heatid="40070" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:31.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.68" eventid="1173" heatid="40131" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:59.68" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.71" eventid="1237" heatid="40219" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:25.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fabienne" lastname="Bauer" birthdate="2013-01-01" gender="F" nation="GER" license="450487" athleteid="36906">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.66" eventid="1123" heatid="40033" lane="6">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:00:33.66" />
                </ENTRY>
                <ENTRY entrytime="00:03:16.79" eventid="1143" heatid="40093" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:03:16.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.19" eventid="1207" heatid="40168" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:39.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:32.91" eventid="1227" heatid="40194" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:32.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.82" eventid="1287" heatid="40314" lane="7">
                  <MEETINFO name="Schwimmfest zum Jahrestag der Schwimmhalle" city="Forst" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:37.70" />
                </ENTRY>
                <ENTRY entrytime="00:03:04.53" eventid="1307" heatid="40351" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:03:04.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.95" eventid="1327" heatid="40384" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:28.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Gustav" lastname="Gärtner" birthdate="2006-01-01" gender="M" nation="GER" license="344042" athleteid="36927">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.13" eventid="1133" heatid="40085" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:25.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.81" eventid="1153" heatid="40109" lane="8">
                  <MEETINFO name="14. Sängerpokal" city="Finsterwalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:43.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.69" eventid="1217" heatid="40187" lane="4">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:31.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.08" eventid="1237" heatid="40229" lane="4">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:01:08.08" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Meike" lastname="Rothe" birthdate="2007-01-01" gender="F" nation="GER" license="345240" athleteid="36936">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.67" eventid="1123" heatid="40051" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:29.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.61" eventid="1163" heatid="40125" lane="8">
                  <MEETINFO name="14. Sängerpokal" city="Finsterwalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:37.61" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.12" eventid="1187" heatid="40149" lane="6">
                  <MEETINFO name="14. Sängerpokal" city="Finsterwalde" course="SCM" approved="GER" date="2025-05-10" qualificationtime="00:02:45.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.40" eventid="1207" heatid="40171" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:37.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.98" eventid="1227" heatid="40209" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:13.98" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5820" nation="GER" region="12" clubid="38874" name="MSV Bautzen 04 e.V.">
          <ATHLETES>
            <ATHLETE firstname="Emily" lastname="Hansel" birthdate="2012-01-01" gender="F" nation="GER" license="439083" athleteid="38888">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.19" eventid="1267" heatid="40271" lane="2">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:11.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.58" eventid="1287" heatid="40314" lane="2">
                  <MEETINFO name="Double-Pool-Meeting (50m Bahn)" city="Riesa" course="LCM" approved="GER" date="2025-02-08" qualificationtime="00:00:37.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.15" eventid="1347" heatid="40410" lane="2">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:38.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.52" eventid="1367" heatid="40444" lane="8">
                  <MEETINFO name="Double-Pool-Meeting (25m Bahn)" city="Riesa" course="SCM" approved="GER" date="2025-02-08" qualificationtime="00:00:39.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.21" eventid="1387" heatid="40477" lane="5">
                  <MEETINFO name="Double-Pool-Meeting (25m Bahn)" city="Riesa" course="SCM" approved="GER" date="2025-02-08" qualificationtime="00:01:26.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Nils" lastname="Grohmann" birthdate="2013-01-01" gender="M" nation="GER" license="454623" athleteid="38884">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.75" eventid="1277" heatid="40292" lane="4">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:15.75" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.58" eventid="1357" heatid="40423" lane="4">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:48.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.90" eventid="1377" heatid="40463" lane="7">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:39.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hannah" lastname="Grohmann" birthdate="2010-01-01" gender="F" nation="GER" license="435383" athleteid="38878">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.33" eventid="1267" heatid="40278" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:07.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.65" eventid="1287" heatid="40318" lane="4">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:00:34.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.07" eventid="1347" heatid="40413" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:31.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.67" eventid="1367" heatid="40452" lane="1">
                  <MEETINFO name="Double-Pool-Meeting (25m Bahn)" city="Riesa" course="SCM" approved="GER" date="2025-02-08" qualificationtime="00:00:35.67" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.16" eventid="1387" heatid="40479" lane="5">
                  <MEETINFO name="Double-Pool-Meeting (25m Bahn)" city="Riesa" course="SCM" approved="GER" date="2025-02-08" qualificationtime="00:01:19.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lorelai" lastname="Florian" birthdate="2009-01-01" gender="F" nation="GER" license="397577" athleteid="38875">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.45" eventid="1267" heatid="40274" lane="1">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:01:09.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.95" eventid="1287" heatid="40318" lane="2">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3339" nation="GER" region="12" clubid="37945" name="SC Freital">
          <ATHLETES>
            <ATHLETE firstname="Alia" lastname="Lange" birthdate="2009-01-01" gender="F" nation="GER" license="402584" athleteid="37951">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.23" eventid="1123" heatid="40058" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.51" eventid="1267" heatid="40286" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:57.50" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.07" eventid="1307" heatid="40360" lane="3" />
                <ENTRY entrytime="00:02:05.69" eventid="1347" heatid="40420" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:05.02" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jule" lastname="Jang" birthdate="2011-01-01" gender="F" nation="GER" license="425575" athleteid="37956">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.50" eventid="1123" heatid="40057" lane="4">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:27.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.06" eventid="1207" heatid="40173" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-11" qualificationtime="00:00:34.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.54" eventid="1267" heatid="40286" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:58.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.77" eventid="1307" heatid="40360" lane="5">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:02:30.47" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.03" eventid="1347" heatid="40420" lane="6">
                  <MEETINFO name="Deutsche Jahrgangsmeisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-13" qualificationtime="00:02:09.03" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Luis Max" lastname="Tetzlaff" birthdate="2013-01-01" gender="M" nation="GER" license="445646" athleteid="37962">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.19" eventid="1133" heatid="40072" lane="6">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:30.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.87" eventid="1217" heatid="40179" lane="4">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:39.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.32" eventid="1237" heatid="40224" lane="7">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:01:17.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.67" eventid="1297" heatid="40336" lane="5">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:33.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.90" eventid="1317" heatid="40370" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:41.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.19" eventid="1357" heatid="40428" lane="3">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:02:28.19" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Moritz-Joy" lastname="Schmidt" birthdate="2006-01-01" gender="M" nation="GER" license="347127" athleteid="37946">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.05" eventid="1133" heatid="40088" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:24.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.28" eventid="1217" heatid="40189" lane="1">
                  <MEETINFO name="41. Goslarer Adler Int. Schwimm-Meeting" city="Goslar" course="SCM" approved="GER" date="2025-03-02" qualificationtime="00:00:31.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.90" eventid="1297" heatid="40347" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:25.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.31" eventid="1377" heatid="40473" lane="7">
                  <MEETINFO name="Plauener Herbst- Mehrkampf" city="Plauen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:28.54" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4581" nation="GER" region="02" clubid="34846" name="VSC 1862 Donauwörth">
          <ATHLETES>
            <ATHLETE firstname="Elena" lastname="Hauser" birthdate="2013-01-01" gender="F" nation="GER" license="458548" athleteid="34847">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.55" eventid="1123" heatid="40052" lane="3">
                  <MEETINFO name="20. Internationaler Sprintpokal" city="Kempten" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:29.49" />
                </ENTRY>
                <ENTRY entrytime="00:03:08.10" eventid="1143" heatid="40095" lane="7">
                  <MEETINFO name="16. internationaler Cool Swimming Cup" city="Gersthofen" course="SCM" approved="GER" date="2025-03-08" qualificationtime="00:03:08.10" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.78" eventid="1163" heatid="40126" lane="2">
                  <MEETINFO name="5. Ingolstädter Nachwuchsschwimmfest" city="Ingolstadt" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:02:31.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.94" eventid="1227" heatid="40211" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:10.94" />
                </ENTRY>
                <ENTRY entrytime="00:04:53.92" eventid="1247" heatid="40243" lane="4">
                  <MEETINFO name="Bayerische aquafeel Jahrgangsmeisterschaften" city="Regensburg" course="LCM" approved="GER" date="2025-07-18" qualificationtime="00:04:53.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.86" eventid="1267" heatid="40283" lane="8">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:03.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.93" eventid="1307" heatid="40360" lane="1">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:33.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.17" eventid="1327" heatid="40386" lane="8">
                  <MEETINFO name="20. Internationaler Sprintpokal" city="Kempten" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:24.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.84" eventid="1347" heatid="40419" lane="6">
                  <MEETINFO name="Bayerische aquafeel Kurzbahnmeisterschaften" city="Nürnberg" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:02:16.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.06" eventid="1387" heatid="40483" lane="2">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:01:10.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3354" nation="GER" region="12" clubid="36842" name="SC DHfK Leipzig">
          <ATHLETES>
            <ATHLETE firstname="Luise" lastname="Kirschner" birthdate="2013-01-01" gender="F" nation="GER" license="446727" athleteid="36880">
              <ENTRIES>
                <ENTRY entrytime="00:06:00.00" eventid="1063" heatid="39995" lane="6" />
                <ENTRY entrytime="00:00:34.82" eventid="1123" heatid="40030" lane="2">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:34.82" />
                </ENTRY>
                <ENTRY entrytime="00:03:27.11" eventid="1143" heatid="40091" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:03:27.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.57" eventid="1207" heatid="40160" lane="7">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:44.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.85" eventid="1267" heatid="40265" lane="2">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:17.85" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.74" eventid="1307" heatid="40350" lane="6">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:03:05.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:38.14" eventid="1327" heatid="40380" lane="1">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:38.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Niels" lastname="Hacker" birthdate="2009-01-01" gender="M" nation="GER" license="381491" athleteid="36850">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.87" eventid="1133" heatid="40084" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:25.72" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.74" eventid="1197" heatid="40154" lane="5">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:02:29.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.48" eventid="1237" heatid="40228" lane="2" />
                <ENTRY entrytime="00:00:59.40" eventid="1277" heatid="40307" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:56.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.82" eventid="1317" heatid="40372" lane="4">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:30.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.07" eventid="1397" heatid="40494" lane="8">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:02.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Teresa Nela" lastname="Hartung" birthdate="2011-01-01" gender="F" nation="GER" license="408424" athleteid="36865">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.46" eventid="1123" heatid="40031" lane="3">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:00:34.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:59.35" eventid="1163" heatid="40116" lane="3">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:59.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.52" eventid="1227" heatid="40197" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:23.33" />
                </ENTRY>
                <ENTRY entrytime="00:03:05.00" eventid="1307" heatid="40350" lane="5">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:03:06.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.07" eventid="1347" heatid="40407" lane="1">
                  <MEETINFO name="34. Nachwuchsschwimmfest des Erfurter SSC" city="Erfurt" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:02:50.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.63" eventid="1367" heatid="40443" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:38.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Vincent" lastname="Hartmann" birthdate="2014-01-01" gender="M" nation="GER" license="459949" athleteid="36857">
              <ENTRIES>
                <ENTRY entrytime="00:21:30.00" eventid="1113" heatid="40023" lane="8" />
                <ENTRY entrytime="00:00:34.28" eventid="1133" heatid="40064" lane="2">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:32.38" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.52" eventid="1237" heatid="40217" lane="8">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:20.05" />
                </ENTRY>
                <ENTRY entrytime="00:05:29.44" eventid="1257" heatid="40249" lane="5">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:05:29.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.05" eventid="1277" heatid="40290" lane="6">
                  <MEETINFO name="Finale Kinderpokal Sachsen" city="Plauen" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:11.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.31" eventid="1357" heatid="40425" lane="2">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:37.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.35" eventid="1377" heatid="40463" lane="4">
                  <MEETINFO name="Schwimmfest unterm Tannenbaum" city="Riesa" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:36.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Waizmann" birthdate="2012-01-01" gender="F" nation="GER" license="442586" athleteid="36888">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.11" eventid="1123" heatid="40032" lane="2">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:34.11" />
                </ENTRY>
                <ENTRY entrytime="00:03:30.00" eventid="1143" heatid="40091" lane="7">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-30" qualificationtime="00:03:34.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.00" eventid="1207" heatid="40161" lane="2">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:44.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.00" eventid="1267" heatid="40266" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:18.98" />
                </ENTRY>
                <ENTRY entrytime="00:03:08.55" eventid="1307" heatid="40350" lane="8">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:03:08.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.00" eventid="1327" heatid="40380" lane="6">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:01:39.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mio Moritz" lastname="Milbach" birthdate="2011-01-01" gender="M" nation="GER" license="408265" athleteid="38612">
              <ENTRIES>
                <ENTRY entrytime="00:11:04.90" eventid="1093" heatid="40014" lane="1" />
                <ENTRY entrytime="00:00:30.73" eventid="1133" heatid="40071" lane="5">
                  <MEETINFO name="31. Lipsiade Stadtsportspiele der Stadt Leipzig" city="Leipzig" course="LCM" approved="GER" date="2025-06-14" qualificationtime="00:00:30.73" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.58" eventid="1153" heatid="40106" lane="2">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:03:03.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.41" eventid="1217" heatid="40179" lane="2">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:00:40.41" />
                </ENTRY>
                <ENTRY entrytime="00:05:22.45" eventid="1257" heatid="40251" lane="7">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:05:22.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.15" eventid="1277" heatid="40296" lane="4">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-25" qualificationtime="00:01:09.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.59" eventid="1317" heatid="40370" lane="8">
                  <MEETINFO name="Int. Dresdner Frühjahrspreis" city="Dresden" course="LCM" approved="GER" date="2025-03-29" qualificationtime="00:02:44.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.79" eventid="1377" heatid="40466" lane="4">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:36.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.90" eventid="1397" heatid="40489" lane="7">
                  <MEETINFO name="Mitteldeutsche Meisterschaften" city="Halle (Saale)" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:20.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marleen" lastname="Forner" birthdate="2011-01-01" gender="F" nation="GER" license="426142" athleteid="36843">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.26" eventid="1123" heatid="40038" lane="7">
                  <MEETINFO name="offene Sächsische Landesmeisterschaften" city="Leipzig" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:00:32.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.60" eventid="1163" heatid="40121" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:02:40.13" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.32" eventid="1227" heatid="40204" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:01:15.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.40" eventid="1287" heatid="40319" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:00:34.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.79" eventid="1307" heatid="40353" lane="4">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:02:54.79" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.95" eventid="1387" heatid="40479" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:01:18.78" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fenja" lastname="Junge" birthdate="2006-01-01" gender="F" nation="GER" license="357784" athleteid="36872">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.67" eventid="1123" heatid="40051" lane="5" />
                <ENTRY entrytime="00:02:59.73" eventid="1143" heatid="40097" lane="4" />
                <ENTRY entrytime="00:00:37.26" eventid="1207" heatid="40171" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:38.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.92" eventid="1267" heatid="40281" lane="2">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:01:07.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.89" eventid="1287" heatid="40325" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:33.51" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.74" eventid="1307" heatid="40359" lane="2">
                  <MEETINFO name="15. Leutzscher Löwenpokal" city="Leipzig" course="LCM" approved="GER" date="2025-01-19" qualificationtime="00:02:41.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.34" eventid="1327" heatid="40389" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:22.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3599" nation="GER" region="13" clubid="38461" name="SV Rotation Halle">
          <ATHLETES>
            <ATHLETE firstname="Daniel" lastname="Nedoborovsky" birthdate="2005-01-01" gender="M" nation="GER" license="342084" athleteid="38467">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.32" eventid="1277" heatid="40305" lane="2">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:00.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.95" eventid="1297" heatid="40340" lane="5">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:30.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.38" eventid="1337" heatid="40398" lane="7">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:01:21.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leonard Edgar" lastname="Bork" birthdate="2010-01-01" gender="M" nation="GER" license="438786" athleteid="38462">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.45" eventid="1277" heatid="40307" lane="8">
                  <MEETINFO name="16. offene KBM S-A Jg. 2015/2016; 2011 u. älter" city="Dessau" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:59.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.87" eventid="1297" heatid="40340" lane="4">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:30.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.34" eventid="1377" heatid="40471" lane="6">
                  <MEETINFO name="19. Sprintmeeting" city="Schönebeck" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:31.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.59" eventid="1397" heatid="40491" lane="4">
                  <MEETINFO name="Schwimmfest anlässlich Luthers Hochzeit" city="Wittenberg" course="SCM" approved="GER" date="2025-06-14" qualificationtime="00:01:10.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="0000" nation="POL" clubid="35898" name="Unia Oświęcim">
          <CONTACT city="Oświęcim" email="p.woznicki@myswimming.pl" name="Woźnicki Piotr" phone="+48 501 042 671" state="MAL" street="Chemików" zip="32-600" />
          <ATHLETES>
            <ATHLETE firstname="Szymon" lastname="Tokarski" birthdate="2010-01-01" gender="M" nation="POL" athleteid="35899">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.07" entrycourse="LCM" eventid="1133" heatid="40087" lane="4">
                </ENTRY>
                <ENTRY entrytime="00:00:29.69" entrycourse="LCM" eventid="1217" heatid="40190" lane="8">
                </ENTRY>
                <ENTRY entrytime="00:01:05.96" entrycourse="LCM" eventid="1337" heatid="40403" lane="1">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="7124" nation="GER" region="12" clubid="37827" name="SV Schneeberg Schwimmen">
          <ATHLETES>
            <ATHLETE firstname="Ben" lastname="Güßmann" birthdate="2011-01-01" gender="M" nation="GER" license="425179" athleteid="37828">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.39" eventid="1133" heatid="40081" lane="6">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:26.90" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.24" eventid="1217" heatid="40183" lane="4">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:33.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.40" eventid="1277" heatid="40301" lane="2">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:01:01.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.12" eventid="1297" heatid="40339" lane="4">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:30.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.93" eventid="1337" heatid="40397" lane="2">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:14.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fiona" lastname="Heymann" birthdate="2011-01-01" gender="F" nation="GER" license="425180" athleteid="37834">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.86" eventid="1123" heatid="40041" lane="2">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:31.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.45" eventid="1287" heatid="40315" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:34.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Janne" lastname="Reichel" birthdate="2009-01-01" gender="M" nation="GER" license="411557" athleteid="37841">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.15" eventid="1133" heatid="40079" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:27.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.82" eventid="1277" heatid="40304" lane="6">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:59.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.85" eventid="1297" heatid="40337" lane="4">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:31.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.74" eventid="1377" heatid="40467" lane="8">
                  <MEETINFO name="Finale Kreis-, Kinder- und Jugendspiele Erzgebirge" city="Zschopau" course="SCM" approved="GER" date="2025-06-15" qualificationtime="00:00:34.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lilly" lastname="Naumann" birthdate="2011-01-01" gender="F" nation="GER" license="432056" athleteid="37837">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.95" eventid="1123" heatid="40030" lane="7">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:00:33.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.96" eventid="1207" heatid="40161" lane="6">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:00:42.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.77" eventid="1367" heatid="40443" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:37.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lucia Zoe" lastname="Veith" birthdate="2010-01-01" gender="F" nation="GER" license="477899" athleteid="37856">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.63" eventid="1123" heatid="40036" lane="5">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:31.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:24.72" eventid="1227" heatid="40198" lane="8">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-13" qualificationtime="00:01:20.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.57" eventid="1367" heatid="40445" lane="4">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:36.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Louis" lastname="Rößler" birthdate="2004-01-01" gender="M" nation="GER" license="297284" athleteid="37846">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.96" eventid="1277" heatid="40307" lane="3">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:55.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.17" eventid="1297" heatid="40343" lane="8">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:27.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.70" eventid="1397" heatid="40491" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:01:03.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Uhlig" birthdate="2013-01-01" gender="F" nation="GER" license="451879" athleteid="37850">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.56" eventid="1123" heatid="40043" lane="7">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:30.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.65" eventid="1207" heatid="40165" lane="5">
                  <MEETINFO name="Auer Wismutpokal" city="Aue" course="SCM" approved="GER" date="2025-09-14" qualificationtime="00:00:39.36" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.80" eventid="1267" heatid="40269" lane="1">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:01:09.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.00" eventid="1287" heatid="40314" lane="1">
                  <MEETINFO name="Bezirksjahrgangs- und Bezirksmeisterschaften" city="Zwickau" course="LCM" approved="GER" date="2025-05-10" qualificationtime="00:00:38.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:33.98" eventid="1327" heatid="40381" lane="6">
                  <MEETINFO name="50. IWS – Internationales Weihnachtsschwimmen" city="Kiel" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:01:27.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5993" nation="GER" region="09" clubid="34597" name="Oldenburger SV 1902">
          <ATHLETES>
            <ATHLETE firstname="Luca" lastname="Prunk" birthdate="2007-01-01" gender="M" nation="GER" license="478284" athleteid="34612">
              <ENTRIES>
                <ENTRY entrytime="00:10:00.50" eventid="1093" heatid="40017" lane="1">
                  <MEETINFO name="Internationale Bestenkämpfe - Frühjahrsausgabe" city="Bremen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:10:37.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.77" eventid="1133" heatid="40080" lane="2" />
                <ENTRY entrytime="00:02:48.69" eventid="1173" heatid="40135" lane="1" />
                <ENTRY entrytime="00:01:16.59" eventid="1237" heatid="40224" lane="4" />
                <ENTRY entrytime="00:04:51.49" eventid="1257" heatid="40255" lane="5" />
                <ENTRY entrytime="00:01:01.25" eventid="1277" heatid="40304" lane="8">
                  <MEETINFO name="Internationale Bestenkämpfe - Frühjahrsausgabe" city="Bremen" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:01:03.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.65" eventid="1357" heatid="40431" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Svea" lastname="Güttler" birthdate="2012-01-01" gender="F" nation="GER" license="441247" athleteid="34598">
              <ENTRIES>
                <ENTRY entrytime="00:11:24.16" eventid="1083" heatid="40006" lane="8" />
                <ENTRY entrytime="00:00:30.68" eventid="1123" heatid="40047" lane="6">
                  <MEETINFO name="Bezirks-Kurzbahn- und Bezirksmastersmeistersch." city="Osnabrück" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:30.68" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.26" eventid="1163" heatid="40121" lane="3">
                  <MEETINFO name="Bezirks-Kurzbahn- und Bezirksmastersmeistersch." city="Osnabrück" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:02:45.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.52" eventid="1227" heatid="40205" lane="3">
                  <MEETINFO name="Landesjahrgangsmeisterschaften Kurzbahn" city="Hannover" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:01:16.98" />
                </ENTRY>
                <ENTRY entrytime="00:05:25.72" eventid="1247" heatid="40238" lane="7">
                  <MEETINFO name="Piranha Meeting" city="Hannover" course="LCM" approved="GER" date="2025-02-28" qualificationtime="00:05:25.72" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Hennemann" birthdate="2008-01-01" gender="F" nation="GER" license="399752" athleteid="34603">
              <ENTRIES>
                <ENTRY entrytime="00:10:15.00" eventid="1083" heatid="40010" lane="7" />
                <ENTRY entrytime="00:00:27.54" eventid="1123" heatid="40057" lane="5">
                  <MEETINFO name="BSV-Sprintercup" city="Bremen - Achterdiek" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:00:27.54" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.22" eventid="1187" heatid="40149" lane="2" />
                <ENTRY entrytime="00:05:04.56" eventid="1247" heatid="40242" lane="5">
                  <MEETINFO name="Piranha Meeting" city="Hannover" course="LCM" approved="GER" date="2025-02-28" qualificationtime="00:05:04.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.33" eventid="1267" heatid="40286" lane="8">
                  <MEETINFO name="BSV-Sprintercup" city="Bremen - Achterdiek" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:00.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.17" eventid="1287" heatid="40329" lane="6">
                  <MEETINFO name="Landesmeisterschaften Kurzbahn" city="Hannover" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:29.17" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.74" eventid="1347" heatid="40419" lane="5">
                  <MEETINFO name="Internationale Bestenkämpfe - Frühjahrsausgabe" city="Bremen" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:02:14.74" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.21" eventid="1387" heatid="40485" lane="1">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:01:06.20" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Michael" gender="M" lastname="Schilling" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="6411" nation="GER" region="04" clubid="35092" name="Potsdamer SV">
          <ATHLETES>
            <ATHLETE firstname="Noah" lastname="Schötz" birthdate="2006-01-01" gender="M" nation="GER" license="348583" athleteid="35139">
              <ENTRIES>
                <ENTRY entrytime="00:00:22.93" eventid="1133" heatid="40089" lane="3">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:00:22.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.20" eventid="1237" heatid="40232" lane="2">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:54.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:50.39" eventid="1277" heatid="40311" lane="5">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:00:50.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.61" eventid="1377" heatid="40474" lane="3">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:24.67" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mina" lastname="Weinert" birthdate="2014-01-01" gender="F" nation="GER" license="492960" athleteid="35155">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.71" eventid="1123" heatid="40027" lane="8">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:36.46" />
                </ENTRY>
                <ENTRY entrytime="00:03:25.00" eventid="1163" heatid="40112" lane="5" />
                <ENTRY entrytime="00:01:30.90" eventid="1227" heatid="40194" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:29.45" />
                </ENTRY>
                <ENTRY entrytime="00:03:25.00" eventid="1307" heatid="40349" lane="8" />
                <ENTRY entrytime="00:00:43.04" eventid="1367" heatid="40440" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:39.74" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jan Malte" lastname="Gräfe" birthdate="2007-01-01" gender="M" nation="GER" license="366984" athleteid="35099">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.07" eventid="1153" heatid="40111" lane="4">
                  <MEETINFO name="European Short Course Championships" city="Lublin" course="SCM" approved="GER" date="2025-12-04" qualificationtime="00:02:05.82" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.99" eventid="1217" heatid="40190" lane="5">
                  <MEETINFO name="European Short Course Championships" city="Lublin" course="SCM" approved="GER" date="2025-12-07" qualificationtime="00:00:26.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.32" eventid="1337" heatid="40403" lane="4">
                  <MEETINFO name="European Short Course Championships" city="Lublin" course="SCM" approved="GER" date="2025-12-02" qualificationtime="00:00:57.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.67" eventid="1397" heatid="40497" lane="2">
                  <MEETINFO name="15. Hamburger Sprint Cup" city="Hamburg-Dulsberg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:00:56.67" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Christopher" lastname="Weidner" birthdate="2005-01-01" gender="M" nation="GER" license="316832" athleteid="35149">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.39" eventid="1133" heatid="40089" lane="7">
                  <MEETINFO name="15. Hamburger Sprint Cup" city="Hamburg-Dulsberg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:00:23.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.17" eventid="1217" heatid="40190" lane="6">
                  <MEETINFO name="15. Hamburger Sprint Cup" city="Hamburg-Dulsberg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:28.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.42" eventid="1297" heatid="40347" lane="5">
                  <MEETINFO name="6. OPERA Swim Classics" city="Wuppertal" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:24.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.77" eventid="1337" heatid="40403" lane="3">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:00.77" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.01" eventid="1397" heatid="40497" lane="6">
                  <MEETINFO name="15. Hamburger Sprint Cup" city="Hamburg-Dulsberg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:00:56.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emma Luise" lastname="Schmid" birthdate="2013-01-01" gender="F" nation="GER" license="437007" athleteid="35124">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.54" eventid="1123" heatid="40037" lane="1">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:00:32.36" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.00" eventid="1187" heatid="40148" lane="5">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-12" qualificationtime="00:03:01.05" />
                </ENTRY>
                <ENTRY entrytime="00:05:20.00" eventid="1247" heatid="40239" lane="2">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:05:18.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.98" eventid="1287" heatid="40318" lane="7">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:34.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:52.13" eventid="1307" heatid="40355" lane="6">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:02:48.29" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.00" eventid="1347" heatid="40411" lane="7">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:28.36" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.53" eventid="1387" heatid="40478" lane="3">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:19.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Elise" lastname="Kramke" birthdate="2014-01-01" gender="F" nation="GER" license="443583" athleteid="35110">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.70" eventid="1123" heatid="40047" lane="7">
                  <MEETINFO name="Norddeutscher Nachwuchsländerkampf" city="Berlin" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:30.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.38" eventid="1163" heatid="40123" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:02:34.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.95" eventid="1207" heatid="40165" lane="1">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:00:39.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.71" eventid="1227" heatid="40208" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:12.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.71" eventid="1287" heatid="40324" lane="2">
                  <MEETINFO name="2. Einladungs-/Kaderprüfungswettkampf" city="Potsdam" course="LCM" approved="GER" date="2025-06-28" qualificationtime="00:00:32.42" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.83" eventid="1307" heatid="40357" lane="5">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:39.61" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.07" eventid="1367" heatid="40457" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:32.79" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.95" eventid="1387" heatid="40478" lane="6">
                  <MEETINFO name="Kurzbahnmeisterschaften des LSV Brandenburg e.V." city="Cottbus" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:17.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Aaron" lastname="Leupold" birthdate="2005-01-01" gender="M" nation="GER" license="319394" athleteid="35119">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.12" eventid="1133" heatid="40089" lane="6">
                  <MEETINFO name="6. OPERA Swim Classics" city="Wuppertal" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:22.74" />
                </ENTRY>
                <ENTRY entrytime="00:04:19.79" eventid="1257" heatid="40259" lane="3">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:04:19.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.14" eventid="1277" heatid="40311" lane="3">
                  <MEETINFO name="15. Hamburger Sprint Cup" city="Hamburg-Dulsberg" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:51.14" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.61" eventid="1357" heatid="40438" lane="4">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:54.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Tobias" lastname="Scholz" birthdate="2006-01-01" gender="M" nation="GER" license="352845" athleteid="35132">
              <ENTRIES>
                <ENTRY entrytime="00:04:40.67" eventid="1073" heatid="40002" lane="6">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:04:40.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.10" eventid="1133" heatid="40089" lane="8">
                  <MEETINFO name="Norddeutsche Meisterschaften" city="Hannover" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:00:24.12" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.55" eventid="1197" heatid="40156" lane="4">
                  <MEETINFO name="Nikar-OPEN" city="Heidelberg" course="LCM" approved="GER" date="2025-07-04" qualificationtime="00:02:01.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.95" eventid="1237" heatid="40232" lane="6">
                  <MEETINFO name="6. OPERA Swim Classics" city="Wuppertal" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:57.95" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.17" eventid="1317" heatid="40376" lane="3">
                  <MEETINFO name="15. Hamburger Sprint Cup" city="Hamburg-Dulsberg" course="SCM" approved="GER" date="2025-09-21" qualificationtime="00:02:08.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.12" eventid="1397" heatid="40497" lane="5">
                  <MEETINFO name="29. Offene Landesmeisterschaften" city="Potsdam" course="LCM" approved="GER" date="2025-07-13" qualificationtime="00:00:54.12" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Kenneth" lastname="Bock" birthdate="2006-01-01" gender="M" nation="GER" license="349019" athleteid="35093">
              <ENTRIES>
                <ENTRY entrytime="00:04:45.49" eventid="1073" heatid="40002" lane="1">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:04:45.49" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.59" eventid="1153" heatid="40111" lane="5">
                  <MEETINFO name="European Short Course Championships" city="Lublin" course="SCM" approved="GER" date="2025-12-04" qualificationtime="00:02:04.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.73" eventid="1217" heatid="40190" lane="7">
                  <MEETINFO name="136. Deutsche Meisterschaften im Schwimmen" city="Berlin" course="LCM" approved="GER" date="2025-05-03" qualificationtime="00:00:28.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.25" eventid="1337" heatid="40403" lane="6">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-13" qualificationtime="00:00:59.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.65" eventid="1397" heatid="40497" lane="3">
                  <MEETINFO name="6. OPERA Swim Classics" city="Wuppertal" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:00:55.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Maike Naomi" lastname="Schwarz" birthdate="1994-01-01" gender="F" nation="GER" license="156094" athleteid="35144">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.13" eventid="1123" heatid="40054" lane="5">
                  <MEETINFO name="Nikar-OPEN" city="Heidelberg" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:28.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.52" eventid="1227" heatid="40206" lane="3">
                  <MEETINFO name="Nikar-OPEN" city="Heidelberg" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:17.34" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.60" eventid="1267" heatid="40284" lane="1">
                  <MEETINFO name="Nikar-OPEN" city="Heidelberg" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:01:03.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.82" eventid="1367" heatid="40451" lane="3">
                  <MEETINFO name="Nikar-OPEN" city="Heidelberg" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:35.42" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Melvin" lastname="Imoudu" birthdate="1999-01-01" gender="M" nation="GER" license="228235" athleteid="35104">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.49" eventid="1133" heatid="40089" lane="1">
                  <MEETINFO name="136. Deutsche Meisterschaften im Schwimmen" city="Berlin" course="LCM" approved="GER" date="2025-05-04" qualificationtime="00:00:23.49" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.69" eventid="1153" heatid="40111" lane="6">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:02:11.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.74" eventid="1217" heatid="40190" lane="4">
                  <MEETINFO name="European Short Course Championships" city="Lublin" course="SCM" approved="GER" date="2025-12-06" qualificationtime="00:00:25.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.43" eventid="1337" heatid="40403" lane="5">
                  <MEETINFO name="European Short Course Championships" city="Lublin" course="SCM" approved="GER" date="2025-12-02" qualificationtime="00:00:56.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.96" eventid="1397" heatid="40497" lane="8">
                  <MEETINFO name="Pokalmeeting Alter Fritz" city="Potsdam" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:00:57.96" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Kassander" lastname="Wolf" birthdate="2007-01-01" gender="M" nation="GER" license="342580" athleteid="35161">
              <ENTRIES>
                <ENTRY entrytime="00:04:48.08" eventid="1073" heatid="40001" lane="4" />
                <ENTRY entrytime="00:00:24.71" eventid="1133" heatid="40088" lane="3">
                  <MEETINFO name="16. Offene Kurzbahnmeisterschaften" city="Potsdam" course="SCM" approved="GER" date="2025-10-12" qualificationtime="00:00:24.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.59" eventid="1173" heatid="40142" lane="4">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-14" qualificationtime="00:02:01.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.16" eventid="1237" heatid="40232" lane="5">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:55.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.59" eventid="1297" heatid="40347" lane="8">
                  <MEETINFO name="Berlin Swim Open" city="Berlin" course="LCM" approved="GER" date="2025-04-26" qualificationtime="00:00:26.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.26" eventid="1317" heatid="40376" lane="6">
                  <MEETINFO name="Norddeutsche Meisterschaften" city="Hannover" course="LCM" approved="GER" date="2025-05-17" qualificationtime="00:02:13.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.40" eventid="1377" heatid="40474" lane="5">
                  <MEETINFO name="Deutsche Kurzbahnmeisterschaften" city="Wuppertal" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:00:25.23" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LoTr" nation="CZE" clubid="39075" name="Lokomotiva Trutnov">
          <CONTACT country="CZ" />
          <ATHLETES>
            <ATHLETE firstname="Karolína" lastname="Malíková" birthdate="2003-01-01" gender="F" nation="CZE" athleteid="39076">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.00" eventid="1123" heatid="40058" lane="2" />
                <ENTRY entrytime="00:01:08.00" eventid="1227" heatid="40213" lane="7" />
                <ENTRY entrytime="00:00:37.99" eventid="1207" heatid="40170" lane="3" />
                <ENTRY entrytime="00:01:03.00" eventid="1267" heatid="40283" lane="3" />
                <ENTRY entrytime="00:01:23.00" eventid="1327" heatid="40389" lane="1" />
                <ENTRY entrytime="00:00:32.00" eventid="1367" heatid="40458" lane="4" />
                <ENTRY entrytime="00:00:31.80" eventid="1287" heatid="40326" lane="7" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5680" nation="GER" region="18" clubid="36838" name="SSV Ulm 1846">
          <CONTACT email="ingo.lachnitt@ssvulm1846.de  " />
          <ATHLETES>
            <ATHLETE firstname="Ilja" lastname="Sukhanov" birthdate="2002-01-01" gender="M" nation="GER" license="267403" athleteid="36839">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.50" eventid="1217" heatid="40187" lane="7">
                  <MEETINFO name="Württembergische Masters-Meisterschaften" city="Stuttgart Bad Cannstatt" course="SCM" approved="GER" date="2025-03-16" qualificationtime="00:00:32.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.50" eventid="1297" heatid="40344" lane="8">
                  <MEETINFO name="56. Deutsche Meisterschaft Masters Kurze Strecke" city="Dresden" course="LCM" approved="GER" date="2025-05-30" qualificationtime="00:00:27.33" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ROLL" nation="SUI" region="RSR" clubid="34841" name="Rolle Natation" shortname="Roll">
          <ATHLETES>
            <ATHLETE firstname="Nele Sophie" lastname="Gläser" birthdate="2014-01-20" gender="F" nation="SUI" athleteid="34842">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.90" entrycourse="LCM" eventid="1123" heatid="40050" lane="3">
                </ENTRY>
                <ENTRY entrytime="00:02:42.24" entrycourse="LCM" eventid="1163" heatid="40123" lane="1">
                </ENTRY>
                <ENTRY entrytime="00:01:11.54" entrycourse="LCM" eventid="1227" heatid="40210" lane="5">
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PKLIL" nation="CZE" clubid="35319" name="Plavecky klub Litomysl">
          <CONTACT country="CZ" />
          <ATHLETES>
            <ATHLETE firstname="Sofie" lastname="Štěpánová" birthdate="2014-01-01" gender="F" nation="CZE" athleteid="35321">
              <ENTRIES>
                <ENTRY entrytime="00:11:35.42" eventid="1083" heatid="40004" lane="5" />
                <ENTRY entrytime="00:00:33.21" eventid="1123" heatid="40035" lane="8" />
                <ENTRY entrytime="00:03:04.21" eventid="1163" heatid="40115" lane="2" />
                <ENTRY entrytime="00:01:29.61" eventid="1227" heatid="40195" lane="3" />
                <ENTRY entrytime="00:05:45.21" eventid="1247" heatid="40236" lane="7" />
                <ENTRY entrytime="00:01:14.25" eventid="1267" heatid="40267" lane="4" />
                <ENTRY entrytime="00:00:40.21" eventid="1287" heatid="40312" lane="3" />
                <ENTRY entrytime="00:02:42.61" eventid="1347" heatid="40408" lane="5" />
                <ENTRY entrytime="00:01:32.61" eventid="1387" heatid="40476" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Šplíchal" birthdate="2012-01-01" gender="M" nation="CZE" athleteid="35791">
              <ENTRIES>
                <ENTRY entrytime="00:10:29.69" eventid="1093" heatid="40015" lane="4" />
                <ENTRY entrytime="00:00:31.53" eventid="1133" heatid="40070" lane="8" />
                <ENTRY entrytime="00:03:09.14" eventid="1153" heatid="40105" lane="7" />
                <ENTRY entrytime="00:01:26.42" eventid="1237" heatid="40218" lane="4" />
                <ENTRY entrytime="00:05:08.67" eventid="1257" heatid="40253" lane="6" />
                <ENTRY entrytime="00:00:35.22" eventid="1297" heatid="40335" lane="6" />
                <ENTRY entrytime="00:02:59.45" eventid="1317" heatid="40365" lane="5" />
                <ENTRY entrytime="00:02:43.64" eventid="1357" heatid="40424" lane="8" />
                <ENTRY entrytime="00:01:28.69" eventid="1397" heatid="40488" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Veronika" lastname="Víchová" birthdate="2015-01-01" gender="F" nation="CZE" athleteid="35801">
              <ENTRIES>
                <ENTRY entrytime="00:12:20.18" eventid="1083" heatid="40003" lane="3" />
                <ENTRY entrytime="00:00:37.17" eventid="1123" heatid="40027" lane="6" />
                <ENTRY entrytime="00:03:03.49" eventid="1163" heatid="40115" lane="3" />
                <ENTRY entrytime="00:01:25.87" eventid="1227" heatid="40196" lane="4" />
                <ENTRY entrytime="00:06:02.13" eventid="1247" heatid="40234" lane="4" />
                <ENTRY entrytime="00:00:42.13" eventid="1287" heatid="40312" lane="2" />
                <ENTRY entrytime="00:01:21.81" eventid="1267" heatid="40262" lane="4" />
                <ENTRY entrytime="00:02:51.58" eventid="1347" heatid="40406" lane="4" />
                <ENTRY entrytime="00:00:40.71" eventid="1367" heatid="40442" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Barbora" lastname="Vokasová" birthdate="2013-01-01" gender="F" nation="CZE" athleteid="35320">
              <ENTRIES>
                <ENTRY entrytime="00:11:08.35" eventid="1083" heatid="40006" lane="3" />
                <ENTRY entrytime="00:00:32.10" eventid="1123" heatid="40039" lane="7" />
                <ENTRY entrytime="00:03:26.21" eventid="1143" heatid="40091" lane="5" />
                <ENTRY entrytime="00:00:41.35" eventid="1207" heatid="40164" lane="6" />
                <ENTRY entrytime="00:05:19.24" eventid="1247" heatid="40239" lane="3" />
                <ENTRY entrytime="00:01:10.24" eventid="1267" heatid="40272" lane="5" />
                <ENTRY entrytime="00:01:29.35" eventid="1327" heatid="40384" lane="8" />
                <ENTRY entrytime="00:02:36.21" eventid="1347" heatid="40411" lane="6" />
                <ENTRY entrytime="00:00:38.21" eventid="1367" heatid="40446" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jáchym" lastname="Votrubec" birthdate="2014-01-01" gender="M" nation="CZE" athleteid="35754">
              <ENTRIES>
                <ENTRY entrytime="00:21:55.00" eventid="1113" heatid="40022" lane="4" />
                <ENTRY entrytime="00:00:34.09" eventid="1133" heatid="40064" lane="3" />
                <ENTRY entrytime="00:05:36.87" eventid="1257" heatid="40248" lane="5" />
                <ENTRY entrytime="00:01:13.58" eventid="1277" heatid="40293" lane="3" />
                <ENTRY entrytime="00:03:01.05" eventid="1317" heatid="40365" lane="1" />
                <ENTRY entrytime="00:02:38.32" eventid="1357" heatid="40425" lane="1" />
                <ENTRY entrytime="00:01:32.43" eventid="1397" heatid="40487" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Agáta" lastname="Votrubcová" birthdate="2012-01-01" gender="F" nation="CZE" athleteid="35762">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.60" eventid="1123" heatid="40047" lane="4" />
                <ENTRY entrytime="00:03:08.94" eventid="1143" heatid="40095" lane="8" />
                <ENTRY entrytime="00:00:38.15" eventid="1207" heatid="40170" lane="8" />
                <ENTRY entrytime="00:05:20.54" eventid="1247" heatid="40239" lane="7" />
                <ENTRY entrytime="00:01:05.70" eventid="1267" heatid="40280" lane="1" />
                <ENTRY entrytime="00:00:32.49" eventid="1287" heatid="40325" lane="8" />
                <ENTRY entrytime="00:01:25.36" eventid="1327" heatid="40387" lane="8" />
                <ENTRY entrytime="00:02:24.33" eventid="1347" heatid="40417" lane="8" />
                <ENTRY entrytime="00:00:36.52" eventid="1367" heatid="40450" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Bulvová" birthdate="2013-01-01" gender="F" nation="CZE" athleteid="35772">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.20" eventid="1123" status="WDR" />
                <ENTRY entrytime="00:03:39.31" eventid="1143" status="WDR" />
                <ENTRY entrytime="00:00:43.39" eventid="1207" status="WDR" />
                <ENTRY entrytime="00:01:33.17" eventid="1227" status="WDR" />
                <ENTRY entrytime="00:01:15.63" eventid="1267" status="WDR" />
                <ENTRY entrytime="00:00:37.46" eventid="1287" status="WDR" />
                <ENTRY entrytime="00:00:41.85" eventid="1367" status="WDR" />
                <ENTRY entrytime="00:01:31.00" eventid="1387" status="WDR" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Eva" lastname="Motyčková " birthdate="2015-01-01" gender="F" nation="CZE" athleteid="35322">
              <ENTRIES>
                <ENTRY entrytime="00:12:19.31" eventid="1083" heatid="40003" lane="5" />
                <ENTRY entrytime="00:00:34.25" eventid="1123" heatid="40032" lane="8" />
                <ENTRY entrytime="00:02:54.69" eventid="1163" heatid="40118" lane="8" />
                <ENTRY entrytime="00:00:44.60" eventid="1207" heatid="40160" lane="1" />
                <ENTRY entrytime="00:01:23.48" eventid="1227" heatid="40199" lane="6" />
                <ENTRY entrytime="00:01:13.94" eventid="1267" heatid="40268" lane="1" />
                <ENTRY entrytime="00:03:00.60" eventid="1307" heatid="40351" lane="4" />
                <ENTRY entrytime="00:00:38.41" eventid="1367" heatid="40446" lane="3" />
                <ENTRY entrytime="00:02:40.23" eventid="1347" heatid="40409" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Adéla" lastname="Štěpánová " birthdate="2015-01-01" gender="F" nation="CZE" athleteid="35323">
              <ENTRIES>
                <ENTRY entrytime="00:12:16.31" eventid="1083" heatid="40003" lane="4" />
                <ENTRY entrytime="00:03:22.13" eventid="1143" heatid="40092" lane="3" />
                <ENTRY entrytime="00:03:07.50" eventid="1163" heatid="40114" lane="3" />
                <ENTRY entrytime="00:01:30.35" eventid="1227" heatid="40195" lane="1" />
                <ENTRY entrytime="00:06:08.23" eventid="1247" heatid="40234" lane="5" />
                <ENTRY entrytime="00:01:13.69" eventid="1267" heatid="40268" lane="3" />
                <ENTRY entrytime="00:02:38.61" eventid="1347" heatid="40410" lane="1" />
                <ENTRY entrytime="00:01:37.21" eventid="1387" heatid="40476" lane="6" />
                <ENTRY entrytime="00:01:35.23" eventid="1327" heatid="40380" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Alena" lastname="Renzová" birthdate="2011-01-01" gender="F" nation="CZE" athleteid="35781">
              <ENTRIES>
                <ENTRY entrytime="00:10:58.42" eventid="1083" heatid="40008" lane="8" />
                <ENTRY entrytime="00:00:33.22" eventid="1123" heatid="40034" lane="4" />
                <ENTRY entrytime="00:03:04.63" eventid="1163" heatid="40115" lane="1" />
                <ENTRY entrytime="00:01:22.98" eventid="1227" heatid="40200" lane="1" />
                <ENTRY entrytime="00:05:14.25" eventid="1247" heatid="40241" lane="7" />
                <ENTRY entrytime="00:01:12.58" eventid="1267" heatid="40270" lane="8" />
                <ENTRY entrytime="00:03:03.90" eventid="1307" heatid="40351" lane="1" />
                <ENTRY entrytime="00:02:41.16" eventid="1347" heatid="40409" lane="2" />
                <ENTRY entrytime="00:00:38.75" eventid="1367" heatid="40445" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3370" nation="GER" region="12" clubid="36302" name="SSV Freiberg">
          <ATHLETES>
            <ATHLETE firstname="Merten" lastname="Kottowski" birthdate="2007-01-01" gender="M" nation="GER" license="367626" athleteid="36307">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.16" eventid="1133" heatid="40087" lane="3">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:25.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.66" eventid="1217" heatid="40185" lane="1">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:35.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.80" eventid="1277" heatid="40309" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:00:56.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.76" eventid="1297" heatid="40342" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:29.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hannah" lastname="Kirchhübel" birthdate="2013-01-01" gender="F" nation="GER" license="446897" athleteid="36303">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.54" eventid="1123" heatid="40052" lane="4">
                  <MEETINFO name="71. Süddeutscher Jugendländervergleich" city="Frankfurt-Höchst" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:29.17" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.25" eventid="1163" heatid="40122" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:43.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.56" eventid="1227" heatid="40207" lane="5">
                  <MEETINFO name="Plauener Herbst- Mehrkampf" city="Plauen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:12.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ingrid" lastname="Lampke" birthdate="2012-01-01" gender="F" nation="GER" license="433827" athleteid="36312">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.17" eventid="1123" heatid="40054" lane="3">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:00:28.20" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.05" eventid="1207" heatid="40164" lane="4">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-30" qualificationtime="00:00:40.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.69" eventid="1267" heatid="40280" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:01:01.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Fynn Luca" lastname="Orosz" birthdate="2007-01-01" gender="M" nation="GER" license="370206" athleteid="36316">
              <ENTRIES>
                <ENTRY entrytime="00:02:35.81" eventid="1153" heatid="40110" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:02:25.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.92" eventid="1217" heatid="40189" lane="6">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:30.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.13" eventid="1297" heatid="40345" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-31" qualificationtime="00:00:26.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.57" eventid="1337" heatid="40402" lane="6">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-29" qualificationtime="00:01:04.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.98" eventid="1397" heatid="40495" lane="4">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:00:58.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Terasa" birthdate="2007-01-01" gender="M" nation="GER" license="363737" athleteid="36328">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.57" eventid="1277" heatid="40309" lane="7">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-06-01" qualificationtime="00:00:54.76" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.50" eventid="1297" heatid="40345" lane="2">
                  <MEETINFO name="Plauener Herbst- Mehrkampf" city="Plauen" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:26.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.00" eventid="1357" heatid="40435" lane="1">
                  <MEETINFO name="26rd Danish International Swim Cup" city="Esbjerg" course="SCM" approved="GER" date="2025-05-30" qualificationtime="00:02:04.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Florentine" lastname="Schmidt" birthdate="2011-01-01" gender="F" nation="GER" license="419436" athleteid="36322">
              <ENTRIES>
                <ENTRY entrytime="00:20:03.55" eventid="1103" heatid="40021" lane="2" />
                <ENTRY entrytime="00:00:29.75" eventid="1123" heatid="40051" lane="7">
                  <MEETINFO name="32. Adventsschwimmfest Erfurt" city="Erfurt" course="LCM" approved="GER" date="2025-11-29" qualificationtime="00:00:29.73" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.96" eventid="1163" heatid="40124" lane="3">
                  <MEETINFO name="Bezirksjahrgangs- und Bezirksmeisterschaften" city="Chemnitz" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:02:29.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.78" eventid="1227" heatid="40207" lane="3">
                  <MEETINFO name="Bezirksjahrgangs- und Bezirksmeisterschaften" city="Chemnitz" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:09.67" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.45" eventid="1267" heatid="40279" lane="7">
                  <MEETINFO name="Bezirksjahrgangs- und Bezirksmeisterschaften" city="Chemnitz" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:04.12" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3355" nation="GER" region="12" clubid="38866" name="SC Poseidon Radebeul">
          <ATHLETES>
            <ATHLETE firstname="Vincent" lastname="Kätzel" birthdate="2011-01-01" gender="M" nation="GER" license="426562" athleteid="38867">
              <ENTRIES>
                <ENTRY entrytime="00:03:05.83" eventid="1153" heatid="40106" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:03:05.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.35" eventid="1173" heatid="40137" lane="7">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:02:40.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.37" eventid="1297" heatid="40338" lane="2">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.37" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.45" eventid="1317" heatid="40371" lane="8">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-18" qualificationtime="00:02:40.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.62" eventid="1357" heatid="40427" lane="3">
                  <MEETINFO name="15. Internationales Silbererz Swim Meeting" city="Freiberg" course="SCM" approved="GER" date="2025-05-17" qualificationtime="00:02:31.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.15" eventid="1377" heatid="40467" lane="5">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:35.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="40498" name="Kometa Brno">
          <ATHLETES>
            <ATHLETE firstname="Daniel" lastname="Gracik" birthdate="2004-01-01" gender="M" nation="CZE" athleteid="40499">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.48" eventid="1297" heatid="40347" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3240" nation="GER" region="16" clubid="38107" name="Eisenacher SSV">
          <ATHLETES>
            <ATHLETE firstname="Leonhard" lastname="Rose" birthdate="2006-01-01" gender="M" nation="GER" license="362415" athleteid="38137">
              <ENTRIES>
                <ENTRY entrytime="00:04:53.02" eventid="1257" heatid="40255" lane="6">
                  <MEETINFO name="Offene Thüringer Meisterschaften lange Strecke" city="Gera" course="LCM" approved="GER" date="2025-02-15" qualificationtime="00:04:59.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.92" eventid="1277" heatid="40303" lane="4">
                  <MEETINFO name="18. Frühjahrsschwimmfest" city="Wetzlar" course="LCM" approved="GER" date="2025-03-08" qualificationtime="00:01:05.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.35" eventid="1357" heatid="40431" lane="4">
                  <MEETINFO name="18. Frühjahrsschwimmfest" city="Wetzlar" course="LCM" approved="GER" date="2025-03-09" qualificationtime="00:02:25.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Henriette" lastname="Penz" birthdate="2010-01-01" gender="F" nation="GER" license="417844" athleteid="38127">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.14" eventid="1123" heatid="40049" lane="4">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:30.07" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.92" eventid="1227" heatid="40205" lane="2">
                  <MEETINFO name="Herbstschwimmfest, ehemals Einladungsschwimmfest" city="Eisenach" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:17.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.71" eventid="1287" heatid="40318" lane="5">
                  <MEETINFO name="Offenes Thüringer Schwimmertreffen" city="Jena" course="LCM" approved="GER" date="2025-05-10" qualificationtime="00:00:34.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.41" eventid="1347" heatid="40414" lane="5">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:25.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Caroline" lastname="Penz" birthdate="2011-01-01" gender="F" nation="GER" license="417079" athleteid="38122">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.41" eventid="1123" heatid="40053" lane="2">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:29.43" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.92" eventid="1227" heatid="40210" lane="8">
                  <MEETINFO name="Offene Thüringer Meisterschaften" city="Erfurt" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:12.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.22" eventid="1287" heatid="40325" lane="3">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:32.16" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.34" eventid="1367" heatid="40458" lane="2">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:32.26" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Steinbach" birthdate="2012-01-01" gender="F" nation="GER" license="481095" athleteid="38112">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.92" eventid="1123" heatid="40035" lane="4">
                  <MEETINFO name="33. Internationale Geraer Stadtmeisterschaften" city="Gera" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:00:32.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.54" eventid="1227" heatid="40195" lane="5">
                  <MEETINFO name="33. Internationale Geraer Stadtmeisterschaften" city="Gera" course="LCM" approved="GER" date="2025-05-18" qualificationtime="00:01:29.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.84" eventid="1287" heatid="40314" lane="5">
                  <MEETINFO name="Offene Thüringer Meisterschaften" city="Erfurt" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:00:36.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.41" eventid="1367" heatid="40444" lane="1">
                  <MEETINFO name="Einladungsschwimmen" city="Eschwege" course="SCM" approved="GER" date="2025-03-22" qualificationtime="00:00:39.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Max" lastname="Rampolt" birthdate="2008-01-01" gender="M" nation="GER" license="370787" athleteid="38117">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.91" eventid="1133" heatid="40086" lane="3">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:00:25.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.54" eventid="1217" heatid="40188" lane="7">
                  <MEETINFO name="Herbstschwimmfest, ehemals Einladungsschwimmfest" city="Eisenach" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:00:33.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.12" eventid="1297" heatid="40346" lane="8">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:27.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.21" eventid="1397" heatid="40495" lane="6">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:01:01.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Stella - Marie" lastname="Dell" birthdate="2009-01-01" gender="F" nation="GER" license="371330" athleteid="38132">
              <ENTRIES>
                <ENTRY entrytime="00:02:40.15" eventid="1163" heatid="40124" lane="8">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-02" qualificationtime="00:02:40.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.14" eventid="1227" heatid="40208" lane="2">
                  <MEETINFO name="Einladungsschwimmen" city="Eschwege" course="SCM" approved="GER" date="2025-03-22" qualificationtime="00:01:15.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.76" eventid="1267" heatid="40276" lane="8">
                  <MEETINFO name="Einladungsschwimmen" city="Eschwege" course="SCM" approved="GER" date="2025-03-22" qualificationtime="00:01:08.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.42" eventid="1367" heatid="40452" lane="5">
                  <MEETINFO name="Einladungsschwimmen" city="Eschwege" course="SCM" approved="GER" date="2025-03-22" qualificationtime="00:00:35.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Baumbach" birthdate="2010-01-01" gender="M" nation="GER" license="413134" athleteid="38108">
              <ENTRIES>
                <ENTRY entrytime="00:02:44.91" eventid="1153" heatid="40109" lane="6">
                  <MEETINFO name="30. Leisslinger Pokal" city="Halle (Saale)" course="LCM" approved="GER" date="2025-05-24" qualificationtime="00:02:43.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.01" eventid="1217" heatid="40187" lane="2">
                  <MEETINFO name="Blacky Cup" city="Erfurt" course="LCM" approved="GER" date="2025-10-26" qualificationtime="00:00:33.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.42" eventid="1337" heatid="40401" lane="5">
                  <MEETINFO name="Thüringer Kurzbahn-Meisterschaften" city="Gotha" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:13.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4452" nation="GER" region="02" clubid="35744" name="TSV Hohenbrunn-Riemerl.">
          <ATHLETES>
            <ATHLETE firstname="Lilly" lastname="Zöckler" birthdate="2008-01-01" gender="F" nation="GER" license="414291" athleteid="35745">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.62" eventid="1123" heatid="40043" lane="1">
                  <MEETINFO name="DMS – BSV Bezirksdurchgang Oberbayern" city="Holzkirchen" course="SCM" approved="GER" date="2025-02-15" qualificationtime="00:00:30.51" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.63" eventid="1143" heatid="40097" lane="7">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:03:01.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.43" eventid="1187" heatid="40148" lane="4">
                  <MEETINFO name="Kreis-JG-Meisterschaften Lagen &amp; Lange Strecken" city="Unterschleißheim" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:02:49.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.97" eventid="1207" heatid="40166" lane="4">
                  <MEETINFO name="Int. Riemerlinger Herbstschwimmfest" city="Riemerling" course="SCM" approved="GER" date="2025-10-04" qualificationtime="00:00:38.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.17" eventid="1267" heatid="40275" lane="1">
                  <MEETINFO name="DMS – BSV Bezirksdurchgang Oberbayern" city="Holzkirchen" course="SCM" approved="GER" date="2025-02-15" qualificationtime="00:01:07.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.82" eventid="1287" heatid="40324" lane="1">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-05" qualificationtime="00:00:32.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.14" eventid="1327" heatid="40386" lane="3">
                  <MEETINFO name="Obb. Jahrgangsmeisterschaften" city="Ingolstadt" course="LCM" approved="GER" date="2025-07-06" qualificationtime="00:01:26.14" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.71" eventid="1387" heatid="40482" lane="6">
                  <MEETINFO name="DMS-J Landesentscheid Bayern" city="Ingolstadt" course="SCM" approved="GER" date="2025-11-22" qualificationtime="00:01:13.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5621" nation="GER" region="03" clubid="38398" name="SG Neukölln e.V. Berlin">
          <ATHLETES>
            <ATHLETE firstname="Immanuel" lastname="Wöhlecke" birthdate="2012-01-01" gender="M" nation="GER" license="446980" athleteid="38454">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.05" eventid="1133" heatid="40064" lane="5">
                  <MEETINFO name="Nachwuchs-Sprinttag des SC Wedding 1929 e.V." city="Berlin" course="SCM" approved="GER" date="2025-11-15" qualificationtime="00:00:33.24" />
                </ENTRY>
                <ENTRY entrytime="00:03:08.72" eventid="1153" heatid="40105" lane="2">
                  <MEETINFO name="8. Int. Neukölln Trophy" city="Berlin" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:03:08.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.76" eventid="1217" heatid="40180" lane="5">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:38.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.52" eventid="1297" heatid="40334" lane="3">
                  <MEETINFO name="8. Int. Neukölln Trophy" city="Berlin" course="SCM" approved="GER" date="2025-10-19" qualificationtime="00:00:35.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.71" eventid="1337" heatid="40396" lane="4">
                  <MEETINFO name="DMSJ Berlin" city="Berlin" course="SCM" approved="GER" date="2025-10-11" qualificationtime="00:01:25.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Wegner" birthdate="2013-01-01" gender="F" nation="GER" license="462447" athleteid="38444">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.36" eventid="1123" heatid="40037" lane="5">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:31.84" />
                </ENTRY>
                <ENTRY entrytime="00:05:38.07" eventid="1247" heatid="40236" lane="4">
                  <MEETINFO name="DMS Landesliga Berlin" city="Berlin" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:05:38.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.71" eventid="1287" heatid="40312" lane="4">
                  <MEETINFO name="Int. Swim-Cup" city="Berlin" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:34.96" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.22" eventid="1347" heatid="40407" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Körsten" birthdate="2012-01-01" gender="F" nation="GER" license="449662" athleteid="38411">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.46" eventid="1123" heatid="40044" lane="8">
                  <MEETINFO name="26. Int. Berolina Cup" city="Berlin" course="LCM" approved="GER" date="2025-02-22" qualificationtime="00:00:31.46" />
                </ENTRY>
                <ENTRY entrytime="00:03:13.74" eventid="1187" heatid="40147" lane="4">
                  <MEETINFO name="DMS Landesliga Berlin" city="Berlin" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:03:15.33" />
                </ENTRY>
                <ENTRY entrytime="00:05:28.00" eventid="1247" heatid="40238" lane="8">
                  <MEETINFO name="25. Int. Wasra-Cup" city="Berlin" course="LCM" approved="GER" date="2025-03-14" qualificationtime="00:05:37.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.31" eventid="1287" heatid="40317" lane="6">
                  <MEETINFO name="Int. Swim-Cup" city="Berlin" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:33.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.22" eventid="1347" heatid="40413" lane="8">
                  <MEETINFO name="25. Int. Wasra-Cup" city="Berlin" course="LCM" approved="GER" date="2025-03-16" qualificationtime="00:02:33.22" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.82" eventid="1387" heatid="40478" lane="4">
                  <MEETINFO name="Int. Swim-Cup" city="Berlin" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:19.27" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Leandra Marie" lastname="Volkmann" birthdate="2003-01-01" gender="F" nation="GER" license="278726" athleteid="38438">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.83" eventid="1123" heatid="40057" lane="2">
                  <MEETINFO name="Offene Berliner Kurzbahnmeisterschaften Masters" city="Berlin" course="SCM" approved="GER" date="2025-11-16" qualificationtime="00:00:28.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.77" eventid="1227" heatid="40213" lane="6">
                  <MEETINFO name="25. Int. Wasra-Cup" city="Berlin" course="LCM" approved="GER" date="2025-03-15" qualificationtime="00:01:07.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.46" eventid="1267" heatid="40285" lane="2">
                  <MEETINFO name="44. Int. Bergbad-Pokal-Schwimmfest" city="Bückeburg" course="LCM" approved="GER" date="2025-06-22" qualificationtime="00:01:02.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.82" eventid="1287" heatid="40326" lane="1">
                  <MEETINFO name="44. Int. Bergbad-Pokal-Schwimmfest" city="Bückeburg" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:00:33.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.67" eventid="1367" heatid="40459" lane="3">
                  <MEETINFO name="28. DMSM Bundesentscheid" city="Nürnberg" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:30.03" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Anne Carola" lastname="Schulz" birthdate="2013-01-01" gender="F" nation="GER" license="435432" athleteid="38425">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.57" eventid="1123" heatid="40048" lane="1">
                  <MEETINFO name="Berliner (Jahrgangs-)Meisterschaften" city="Berlin" course="LCM" approved="GER" date="2025-06-28" qualificationtime="00:00:30.57" />
                </ENTRY>
                <ENTRY entrytime="00:02:57.65" eventid="1163" heatid="40117" lane="8" />
                <ENTRY entrytime="00:05:09.99" eventid="1247" heatid="40242" lane="7">
                  <MEETINFO name="DM Schwimmerischer Mehrkampf" city="Dortmund" course="LCM" approved="GER" date="2025-06-06" qualificationtime="00:05:09.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.09" eventid="1267" heatid="40279" lane="6">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:04.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.82" eventid="1347" heatid="40416" lane="8">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:21.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Schnabel" birthdate="2013-01-01" gender="F" nation="GER" license="475926" athleteid="38418">
              <ENTRIES>
                <ENTRY entrytime="00:03:26.06" eventid="1143" heatid="40091" lane="4">
                  <MEETINFO name="DMS Landesliga Berlin" city="Berlin" course="SCM" approved="GER" date="2025-11-30" qualificationtime="00:03:12.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.99" eventid="1207" heatid="40163" lane="1">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:40.16" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.77" eventid="1267" heatid="40268" lane="7">
                  <MEETINFO name="Int. Swim-Cup" city="Berlin" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:01:13.77" />
                </ENTRY>
                <ENTRY entrytime="00:03:03.56" eventid="1307" heatid="40351" lane="7">
                  <MEETINFO name="Int. Swim-Cup" city="Berlin" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:03:03.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:31.85" eventid="1327" heatid="40382" lane="2">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:01:28.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.67" eventid="1347" heatid="40406" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ronja" lastname="Brandt" birthdate="2010-01-01" gender="F" nation="GER" license="418440" athleteid="38399">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.33" eventid="1123" heatid="40044" lane="6">
                  <MEETINFO name="28. Internationaler Sportbadpokal" city="Berlin" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:00:31.33" />
                </ENTRY>
                <ENTRY entrytime="00:02:53.20" eventid="1143" heatid="40098" lane="5">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-07" qualificationtime="00:02:53.20" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.28" eventid="1207" heatid="40171" lane="5">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:37.28" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.92" eventid="1307" heatid="40359" lane="7">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:02:37.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:22.55" eventid="1327" heatid="40389" lane="2">
                  <MEETINFO name="Int. Swim-Cup" city="Berlin" course="SCM" approved="GER" date="2025-09-28" qualificationtime="00:01:22.55" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Piloka Marie" lastname="Weisner" birthdate="2013-01-01" gender="F" nation="GER" license="472213" athleteid="38449">
              <ENTRIES>
                <ENTRY entrytime="00:01:16.24" eventid="1227" heatid="40206" lane="5">
                  <MEETINFO name="8. Int. Neukölln Trophy" city="Berlin" course="SCM" approved="GER" date="2025-10-18" qualificationtime="00:01:12.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.01" eventid="1267" heatid="40281" lane="1">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:02.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.60" eventid="1287" heatid="40326" lane="5">
                  <MEETINFO name="26. Int. Berolina Cup" city="Berlin" course="LCM" approved="GER" date="2025-02-23" qualificationtime="00:00:31.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.02" eventid="1367" heatid="40453" lane="3">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:00:32.77" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Wilma" lastname="Gottschlich" birthdate="2009-01-01" gender="F" nation="GER" license="389257" athleteid="38405">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.71" eventid="1123" heatid="40055" lane="2">
                  <MEETINFO name="26. Int. Berolina Cup" city="Berlin" course="LCM" approved="GER" date="2025-02-22" qualificationtime="00:00:28.98" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.82" eventid="1227" heatid="40210" lane="1" />
                <ENTRY entrytime="00:01:03.78" eventid="1267" heatid="40283" lane="1" />
                <ENTRY entrytime="00:00:32.49" eventid="1287" heatid="40325" lane="1">
                  <MEETINFO name="Int. Swim-Cup" city="Berlin" course="SCM" approved="GER" date="2025-09-27" qualificationtime="00:00:32.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.10" eventid="1367" heatid="40457" lane="2">
                  <MEETINFO name="26. Int. Berolina Cup" city="Berlin" course="LCM" approved="GER" date="2025-02-23" qualificationtime="00:00:33.62" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Noa" lastname="Ulucay" birthdate="2012-01-01" gender="M" nation="GER" license="456363" athleteid="38431">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.84" eventid="1133" heatid="40069" lane="2">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-09" qualificationtime="00:00:29.46" />
                </ENTRY>
                <ENTRY entrytime="00:03:02.45" eventid="1173" heatid="40131" lane="8" />
                <ENTRY entrytime="00:01:24.01" eventid="1237" heatid="40219" lane="4">
                  <MEETINFO name="44. Int. Bergbad-Pokal-Schwimmfest" city="Bückeburg" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:01:24.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.45" eventid="1277" heatid="40295" lane="8">
                  <MEETINFO name="Berliner Kurzbahnmeisterschaften" city="Berlin" course="SCM" approved="GER" date="2025-11-08" qualificationtime="00:01:05.18" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.84" eventid="1357" heatid="40426" lane="3">
                  <MEETINFO name="28. Internationaler Sportbadpokal" city="Berlin" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:02:34.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.13" eventid="1397" heatid="40488" lane="5">
                  <MEETINFO name="28. Internationaler Sportbadpokal" city="Berlin" course="LCM" approved="GER" date="2025-06-07" qualificationtime="00:01:25.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.34" eventid="1183" heatid="40144" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="38438" number="1" />
                    <RELAYPOSITION athleteid="38399" number="2" />
                    <RELAYPOSITION athleteid="38405" number="3" />
                    <RELAYPOSITION athleteid="38449" number="4" />
                  </RELAYPOSITIONS>
                  <MEETINFO name="8. Int. Neukölln Trophy" city="Berlin" date="2025-10-19" qualificationtime="00:02:08.46" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="3337" nation="GER" region="12" clubid="38928" name="SV Lok Görlitz e.V.">
          <ATHLETES>
            <ATHLETE firstname="Nelly" lastname="Eifler" birthdate="2014-01-01" gender="F" nation="GER" license="451392" athleteid="38938">
              <ENTRIES>
                <ENTRY entrytime="00:01:17.80" eventid="1267" heatid="40265" lane="6">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:17.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.62" eventid="1287" heatid="40317" lane="1">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:35.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.99" eventid="1367" heatid="40444" lane="4">
                  <MEETINFO name="Bezirks-Kurzbahnmeistersch. JG 2016 u.ä." city="Riesa" course="SCM" approved="GER" date="2025-09-20" qualificationtime="00:00:37.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marah" lastname="Tschirner" birthdate="2012-01-01" gender="F" nation="GER" license="442928" athleteid="38965">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.14" eventid="1267" heatid="40268" lane="8">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-12" qualificationtime="00:01:14.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.88" eventid="1287" heatid="40316" lane="5">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:34.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.56" eventid="1367" heatid="40446" lane="8">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:37.83" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Vincent" lastname="Steudtner" birthdate="2012-01-01" gender="M" nation="GER" license="442934" athleteid="38960">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.13" eventid="1133" heatid="40082" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:26.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.11" eventid="1237" heatid="40228" lane="3">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:06.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.37" eventid="1277" heatid="40305" lane="1">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:00:58.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.39" eventid="1297" heatid="40341" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:29.20" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Aurelius" lastname="Vogt" birthdate="2013-01-01" gender="M" nation="GER" license="445775" athleteid="38973">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.99" eventid="1133" heatid="40076" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:28.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.09" eventid="1173" heatid="40135" lane="2">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:42.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.27" eventid="1237" heatid="40225" lane="1">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:11.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.13" eventid="1277" heatid="40299" lane="6">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:04.28" />
                </ENTRY>
                <ENTRY entrytime="00:02:47.41" eventid="1317" heatid="40369" lane="1">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:40.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.64" eventid="1377" heatid="40469" lane="6">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:32.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Pepe" lastname="Tzschoppe" birthdate="2011-01-01" gender="M" nation="GER" license="400384" athleteid="38969">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.81" eventid="1133" heatid="40080" lane="7">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:00:27.81" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.11" eventid="1173" heatid="40138" lane="3">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:28.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.12" eventid="1237" heatid="40227" lane="5">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:08.46" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Louis Matthias" lastname="Dietrich" birthdate="2011-01-01" gender="M" nation="GER" license="425561" athleteid="38933">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.93" eventid="1133" heatid="40079" lane="4">
                  <MEETINFO name="Kreis-Kinder- und Jugendspiele Jg. 2015 - 2007" city="Görlitz" course="SCM" approved="GER" date="2025-05-24" qualificationtime="00:00:27.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.11" eventid="1217" heatid="40184" lane="1">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:33.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.78" eventid="1297" heatid="40339" lane="6">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:30.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.11" eventid="1337" heatid="40398" lane="2">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:01:17.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jette" lastname="Gunsilius" birthdate="2011-01-01" gender="F" nation="GER" license="425560" athleteid="38942">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.16" eventid="1267" heatid="40278" lane="4">
                  <MEETINFO name="27. Schwimmfest am Windberg" city="Freital" course="SCM" approved="GER" date="2025-06-28" qualificationtime="00:01:05.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.53" eventid="1307" heatid="40355" lane="4">
                  <MEETINFO name="6. Mehrkampfwettkampf" city="Berlin-Marzahn" course="LCM" approved="GER" date="2025-04-05" qualificationtime="00:02:50.53" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.79" eventid="1347" heatid="40413" lane="2">
                  <MEETINFO name="Bezirksmeisterschaften der Jahrgänge 2017 u.ä." city="Dresden" course="LCM" approved="GER" date="2025-04-13" qualificationtime="00:02:30.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Julian" lastname="Bormann" birthdate="2012-01-01" gender="M" nation="GER" license="442932" athleteid="38929">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.59" eventid="1133" heatid="40067" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-26" qualificationtime="00:00:30.13" />
                </ENTRY>
                <ENTRY entrytime="00:03:18.11" eventid="1153" heatid="40104" lane="8">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:03:12.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.11" eventid="1217" heatid="40180" lane="7">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:00:37.45" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lynn Xenia" lastname="Illing" birthdate="2012-01-01" gender="F" nation="GER" license="436674" athleteid="38946">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.44" eventid="1123" heatid="40053" lane="8">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:29.44" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.73" eventid="1163" heatid="40123" lane="7">
                  <MEETINFO name="Sparkassen Landesjugendspiele" city="Dresden" course="LCM" approved="GER" date="2025-06-21" qualificationtime="00:02:45.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.24" eventid="1207" heatid="40169" lane="4">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:38.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.79" eventid="1227" heatid="40209" lane="5">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:13.79" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.45" eventid="1267" heatid="40280" lane="3">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:05.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.09" eventid="1287" heatid="40325" lane="5">
                  <MEETINFO name="32. Görlitzer Sprintmeeting" city="Görlitz" course="SCM" approved="GER" date="2025-09-06" qualificationtime="00:00:32.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.43" eventid="1327" heatid="40388" lane="5">
                  <MEETINFO name="offene Sächsische Kurzbahnmeisterschaften" city="Riesa" course="SCM" approved="GER" date="2025-10-25" qualificationtime="00:01:23.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.93" eventid="1367" heatid="40456" lane="8">
                  <MEETINFO name="Kreis-Kinder- und Jugendspiele Jg. 2015 - 2007" city="Görlitz" course="SCM" approved="GER" date="2025-05-24" qualificationtime="00:00:33.93" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lukas" lastname="Nowotny" birthdate="2013-01-01" gender="M" nation="GER" license="445777" athleteid="38955">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.94" eventid="1277" heatid="40292" lane="2">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:10.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:39.46" eventid="1297" heatid="40332" lane="5">
                  <MEETINFO name="Talentewettkampf" city="Cottbus" course="SCM" approved="GER" date="2025-06-22" qualificationtime="00:00:39.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.38" eventid="1337" heatid="40393" lane="6">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:01:32.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.11" eventid="1357" heatid="40424" lane="7">
                  <MEETINFO name="11. Internationaler NEISSE – POKAL" city="Görlitz" course="SCM" approved="GER" date="2025-11-01" qualificationtime="00:02:36.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Wacha" birthdate="2014-01-01" gender="F" nation="GER" license="451399" athleteid="38980">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="1267" heatid="40263" lane="5">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:01:20.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.50" eventid="1287" heatid="40313" lane="5">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:38.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.00" eventid="1367" heatid="40442" lane="1">
                  <MEETINFO name="Herbstschwimmfest des Schwimmbezirk Dresden" city="Dresden" course="LCM" approved="GER" date="2025-11-02" qualificationtime="00:00:41.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="33676" course="LCM" gender="M" name="2007 und älter" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="18" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:12.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:15.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:25.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:15.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33677" course="LCM" gender="F" name="2007 und älter" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="18" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:28.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:45.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33680" course="LCM" gender="M" name="2008" type="MAXIMUM">
      <AGEGROUP agemax="17" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:12.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:25.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:30.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33681" course="LCM" gender="F" name="2008" type="MAXIMUM">
      <AGEGROUP agemax="17" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:15.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:28.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:15.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33678" course="LCM" gender="M" name="2009" type="MAXIMUM">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:12.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:45.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:25.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:45.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33679" course="LCM" gender="F" name="2009" type="MAXIMUM">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:30.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:28.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:45.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33682" course="LCM" gender="M" name="2010" type="MAXIMUM">
      <AGEGROUP agemax="15" agemin="15" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:18.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:25.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:09.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:15.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33683" course="LCM" gender="F" name="2010" type="MAXIMUM">
      <AGEGROUP agemax="15" agemin="15" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:41.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:45.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:28.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:15.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33684" course="LCM" gender="M" name="2011" type="MAXIMUM">
      <AGEGROUP agemax="14" agemin="14" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:15.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:50.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:35.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:12.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:45.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33685" course="LCM" gender="F" name="2011" type="MAXIMUM">
      <AGEGROUP agemax="14" agemin="14" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:25.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:00.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:31.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:45.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33686" course="LCM" gender="M" name="2012" type="MAXIMUM">
      <AGEGROUP agemax="13" agemin="13" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:30.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:41.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:30.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:10.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:32.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:50.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:15.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33687" course="LCM" gender="F" name="2012" type="MAXIMUM">
      <AGEGROUP agemax="13" agemin="13" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:35.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:43.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:15.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:36.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:50.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:16.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:15.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33688" course="LCM" gender="M" name="2013" type="MAXIMUM">
      <AGEGROUP agemax="12" agemin="12" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:45.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:44.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:45.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:10.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:35.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:41.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:00.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33689" course="LCM" gender="F" name="2013" type="MAXIMUM">
      <AGEGROUP agemax="12" agemin="12" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:45.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:44.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:30.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:10.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:35.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:41.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:45.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33690" course="LCM" gender="M" name="2014" type="MAXIMUM">
      <AGEGROUP agemax="11" agemin="11" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:47.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:47.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:25.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:15.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:55.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:43.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:20.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:23.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:25.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:44.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:22:00.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33691" course="LCM" gender="F" name="2014" type="MAXIMUM">
      <AGEGROUP agemax="11" agemin="11" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:47.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:47.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:25.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:45.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:55.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:43.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:20.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:23.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:25.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:44.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:22:15.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33692" course="LCM" gender="M" name="2015" type="MAXIMUM">
      <AGEGROUP agemax="10" agemin="10" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:50.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:49.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:00.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:26.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:46.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:41.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:22:45.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="33693" course="LCM" gender="F" name="2015" type="MAXIMUM">
      <AGEGROUP agemax="10" agemin="10" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:50.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:50.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:49.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:30.99">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.99">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:26.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.99">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:46.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:41.99">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:23:30.99">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.99">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>