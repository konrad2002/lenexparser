<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.24" registration="">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Marienberg" course="SCM" name="26. Internationaler Erzgebirgs-Schwimmcup 2023" nation="GER" organizer="Schwimm-Team Erzgebirge e.V." hostclub="Schwimm-Team Erzgebirge e.V." deadline="2023-11-28" timing="AUTOMATIC">
      <CONTACT city="Olbernhau" email="alex@schwimmteamerzgebirge.de" internet="www.schwimmteamerzgebirge.de" name="Steiner, Alexander" phone="+49 373607 5177" street="Hammergasse 24" zip="09526" />
      <AGEDATE type="YEAR" value="2023-01-01" />
      <SESSIONS>
        <SESSION number="1" date="2023-12-09" daytime="08:45" officialmeeting="08:15" warmupfrom="07:30">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="1001" number="1" />
                <HEAT heatid="1002" number="2" />
                <HEAT heatid="1003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="1489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="5" resultid="240" />
                    <RANKING place="2" resultid="590" />
                    <RANKING place="1" resultid="840" />
                    <RANKING place="4" resultid="1354" />
                    <RANKING place="3" resultid="1520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="158" />
                    <RANKING place="2" resultid="290" />
                    <RANKING place="1" resultid="547" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="2" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="2000" number="0" />
                <HEAT heatid="2001" number="1" />
                <HEAT heatid="2002" number="2" />
                <HEAT heatid="2003" number="3" />
                <HEAT heatid="2004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="298" />
                    <RANKING place="1" resultid="1442" />
                    <RANKING place="3" resultid="1448" />
                    <RANKING place="2" resultid="1454" />
                    <RANKING place="5" resultid="1538" />
                    <RANKING place="6" resultid="1815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="8" />
                    <RANKING place="3" resultid="305" />
                    <RANKING place="2" resultid="696" />
                    <RANKING place="4" resultid="1568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="1658" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="3" gender="F" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="3000" number="0" />
                <HEAT heatid="3001" number="1" />
                <HEAT heatid="3002" number="2" />
                <HEAT heatid="3003" number="3" />
                <HEAT heatid="3004" number="4" />
                <HEAT heatid="3005" number="5" />
                <HEAT heatid="3006" number="6" />
                <HEAT heatid="3007" number="7" />
                <HEAT heatid="3008" number="8" />
                <HEAT heatid="3009" number="9" />
                <HEAT heatid="3010" number="10" />
                <HEAT heatid="3011" number="11" />
                <HEAT heatid="3012" number="12" />
                <HEAT heatid="3013" number="13" />
                <HEAT heatid="3014" number="14" />
                <HEAT heatid="3015" number="15" />
                <HEAT heatid="3016" number="16" />
                <HEAT heatid="3017" number="17" />
                <HEAT heatid="3018" number="18" />
                <HEAT heatid="3019" number="19" />
                <HEAT heatid="3020" number="20" />
                <HEAT heatid="3021" number="21" />
                <HEAT heatid="3022" number="22" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="5" resultid="302" />
                    <RANKING place="6" resultid="501" />
                    <RANKING place="4" resultid="575" />
                    <RANKING place="11" resultid="628" />
                    <RANKING place="1" resultid="639" />
                    <RANKING place="10" resultid="645" />
                    <RANKING place="2" resultid="789" />
                    <RANKING place="3" resultid="800" />
                    <RANKING place="7" resultid="858" />
                    <RANKING place="8" resultid="1593" />
                    <RANKING place="12" resultid="1608" />
                    <RANKING place="9" resultid="1750" />
                    <RANKING place="13" resultid="1805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="355" />
                    <RANKING place="8" resultid="516" />
                    <RANKING place="5" resultid="520" />
                    <RANKING place="10" resultid="585" />
                    <RANKING place="7" resultid="685" />
                    <RANKING place="9" resultid="704" />
                    <RANKING place="11" resultid="758" />
                    <RANKING place="4" resultid="954" />
                    <RANKING place="6" resultid="1290" />
                    <RANKING place="3" resultid="1294" />
                    <RANKING place="1" resultid="1298" />
                    <RANKING place="12" resultid="1517" />
                    <RANKING place="13" resultid="1901" />
                    <RANKING place="14" resultid="1926" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="262" />
                    <RANKING place="15" resultid="445" />
                    <RANKING place="9" resultid="691" />
                    <RANKING place="1" resultid="715" />
                    <RANKING place="13" resultid="731" />
                    <RANKING place="7" resultid="747" />
                    <RANKING place="6" resultid="794" />
                    <RANKING place="5" resultid="811" />
                    <RANKING place="2" resultid="935" />
                    <RANKING place="10" resultid="984" />
                    <RANKING place="11" resultid="1153" />
                    <RANKING place="4" resultid="1372" />
                    <RANKING place="14" resultid="1490" />
                    <RANKING place="18" resultid="1532" />
                    <RANKING place="12" resultid="1703" />
                    <RANKING place="17" resultid="1746" />
                    <RANKING place="8" resultid="1800" />
                    <RANKING place="16" resultid="1878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="7" resultid="721" />
                    <RANKING place="14" resultid="770" />
                    <RANKING place="9" resultid="1306" />
                    <RANKING place="4" resultid="1318" />
                    <RANKING place="1" resultid="1325" />
                    <RANKING place="2" resultid="1330" />
                    <RANKING place="11" resultid="1336" />
                    <RANKING place="3" resultid="1342" />
                    <RANKING place="6" resultid="1348" />
                    <RANKING place="10" resultid="1360" />
                    <RANKING place="8" resultid="1521" />
                    <RANKING place="5" resultid="1526" />
                    <RANKING place="12" resultid="1719" />
                    <RANKING place="13" resultid="1763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="10" resultid="35" />
                    <RANKING place="11" resultid="49" />
                    <RANKING place="8" resultid="159" />
                    <RANKING place="16" resultid="319" />
                    <RANKING place="2" resultid="413" />
                    <RANKING place="12" resultid="478" />
                    <RANKING place="3" resultid="525" />
                    <RANKING place="1" resultid="548" />
                    <RANKING place="9" resultid="726" />
                    <RANKING place="4" resultid="1053" />
                    <RANKING place="14" resultid="1145" />
                    <RANKING place="15" resultid="1164" />
                    <RANKING place="19" resultid="1168" />
                    <RANKING place="5" resultid="1366" />
                    <RANKING place="13" resultid="1599" />
                    <RANKING place="7" resultid="1690" />
                    <RANKING place="17" resultid="1789" />
                    <RANKING place="18" resultid="1853" />
                    <RANKING place="6" resultid="1864" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="4" gender="M" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="4000" number="0" />
                <HEAT heatid="4001" number="1" />
                <HEAT heatid="4002" number="2" />
                <HEAT heatid="4003" number="3" />
                <HEAT heatid="4004" number="4" />
                <HEAT heatid="4005" number="5" />
                <HEAT heatid="4006" number="6" />
                <HEAT heatid="4007" number="7" />
                <HEAT heatid="4008" number="8" />
                <HEAT heatid="4009" number="9" />
                <HEAT heatid="4010" number="10" />
                <HEAT heatid="4011" number="11" />
                <HEAT heatid="4012" number="12" />
                <HEAT heatid="4013" number="13" />
                <HEAT heatid="4014" number="14" />
                <HEAT heatid="4015" number="15" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="2" resultid="671" />
                    <RANKING place="1" resultid="1378" />
                    <RANKING place="3" resultid="1895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="6" resultid="236" />
                    <RANKING place="1" resultid="483" />
                    <RANKING place="2" resultid="487" />
                    <RANKING place="3" resultid="491" />
                    <RANKING place="4" resultid="649" />
                    <RANKING place="5" resultid="907" />
                    <RANKING place="7" resultid="990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="554" />
                    <RANKING place="1" resultid="622" />
                    <RANKING place="5" resultid="709" />
                    <RANKING place="8" resultid="885" />
                    <RANKING place="3" resultid="917" />
                    <RANKING place="2" resultid="1436" />
                    <RANKING place="7" resultid="1596" />
                    <RANKING place="10" resultid="1725" />
                    <RANKING place="9" resultid="1729" />
                    <RANKING place="6" resultid="1741" />
                    <RANKING place="11" resultid="1796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="9" resultid="360" />
                    <RANKING place="3" resultid="424" />
                    <RANKING place="1" resultid="697" />
                    <RANKING place="2" resultid="1023" />
                    <RANKING place="5" resultid="1100" />
                    <RANKING place="8" resultid="1390" />
                    <RANKING place="4" resultid="1412" />
                    <RANKING place="7" resultid="1424" />
                    <RANKING place="6" resultid="1430" />
                    <RANKING place="10" resultid="1628" />
                    <RANKING place="11" resultid="1672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="339" />
                    <RANKING place="4" resultid="387" />
                    <RANKING place="1" resultid="531" />
                    <RANKING place="2" resultid="1013" />
                    <RANKING place="3" resultid="1400" />
                    <RANKING place="8" resultid="1550" />
                    <RANKING place="7" resultid="1633" />
                    <RANKING place="5" resultid="1648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="4" resultid="32" />
                    <RANKING place="1" resultid="440" />
                    <RANKING place="5" resultid="542" />
                    <RANKING place="7" resultid="960" />
                    <RANKING place="6" resultid="1048" />
                    <RANKING place="2" resultid="1068" />
                    <RANKING place="3" resultid="1574" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="5" gender="F" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="5000" number="0" />
                <HEAT heatid="5001" number="1" />
                <HEAT heatid="5002" number="2" />
                <HEAT heatid="5003" number="3" />
                <HEAT heatid="5004" number="4" />
                <HEAT heatid="5005" number="5" />
                <HEAT heatid="5006" number="6" />
                <HEAT heatid="5007" number="7" />
                <HEAT heatid="5008" number="8" />
                <HEAT heatid="5009" number="9" />
                <HEAT heatid="5010" number="10" />
                <HEAT heatid="5011" number="11" />
                <HEAT heatid="5012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="5" resultid="537" />
                    <RANKING place="2" resultid="579" />
                    <RANKING place="1" resultid="640" />
                    <RANKING place="4" resultid="801" />
                    <RANKING place="6" resultid="1512" />
                    <RANKING place="7" resultid="1609" />
                    <RANKING place="3" resultid="1751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="5" resultid="517" />
                    <RANKING place="1" resultid="586" />
                    <RANKING place="2" resultid="617" />
                    <RANKING place="3" resultid="686" />
                    <RANKING place="4" resultid="705" />
                    <RANKING place="6" resultid="1902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="692" />
                    <RANKING place="6" resultid="732" />
                    <RANKING place="1" resultid="936" />
                    <RANKING place="5" resultid="1544" />
                    <RANKING place="2" resultid="1605" />
                    <RANKING place="4" resultid="1704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="59" />
                    <RANKING place="3" resultid="274" />
                    <RANKING place="9" resultid="282" />
                    <RANKING place="10" resultid="469" />
                    <RANKING place="11" resultid="771" />
                    <RANKING place="7" resultid="1307" />
                    <RANKING place="12" resultid="1319" />
                    <RANKING place="4" resultid="1349" />
                    <RANKING place="1" resultid="1355" />
                    <RANKING place="5" resultid="1361" />
                    <RANKING place="6" resultid="1527" />
                    <RANKING place="8" resultid="1764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="270" />
                    <RANKING place="11" resultid="320" />
                    <RANKING place="4" resultid="563" />
                    <RANKING place="8" resultid="727" />
                    <RANKING place="1" resultid="1054" />
                    <RANKING place="3" resultid="1131" />
                    <RANKING place="13" resultid="1134" />
                    <RANKING place="10" resultid="1147" />
                    <RANKING place="9" resultid="1600" />
                    <RANKING place="12" resultid="1602" />
                    <RANKING place="5" resultid="1691" />
                    <RANKING place="7" resultid="1755" />
                    <RANKING place="2" resultid="1865" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="6" gender="M" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="6000" number="0" />
                <HEAT heatid="6001" number="1" />
                <HEAT heatid="6002" number="2" />
                <HEAT heatid="6003" number="3" />
                <HEAT heatid="6004" number="4" />
                <HEAT heatid="6005" number="5" />
                <HEAT heatid="6006" number="6" />
                <HEAT heatid="6007" number="7" />
                <HEAT heatid="6008" number="8" />
                <HEAT heatid="6009" number="9" />
                <HEAT heatid="6010" number="10" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="1" resultid="1896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="213" />
                    <RANKING place="1" resultid="1386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="248" />
                    <RANKING place="1" resultid="430" />
                    <RANKING place="5" resultid="710" />
                    <RANKING place="7" resultid="1142" />
                    <RANKING place="6" resultid="1437" />
                    <RANKING place="3" resultid="1455" />
                    <RANKING place="4" resultid="1708" />
                    <RANKING place="8" resultid="1726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="14" />
                    <RANKING place="1" resultid="20" />
                    <RANKING place="3" resultid="306" />
                    <RANKING place="12" resultid="361" />
                    <RANKING place="4" resultid="879" />
                    <RANKING place="10" resultid="1043" />
                    <RANKING place="6" resultid="1413" />
                    <RANKING place="11" resultid="1425" />
                    <RANKING place="7" resultid="1431" />
                    <RANKING place="5" resultid="1569" />
                    <RANKING place="9" resultid="1629" />
                    <RANKING place="8" resultid="1673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="998" />
                    <RANKING place="2" resultid="1095" />
                    <RANKING place="4" resultid="1401" />
                    <RANKING place="6" resultid="1551" />
                    <RANKING place="1" resultid="1590" />
                    <RANKING place="5" resultid="1634" />
                    <RANKING place="7" resultid="1649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="773" />
                    <RANKING place="2" resultid="829" />
                    <RANKING place="4" resultid="1575" />
                    <RANKING place="3" resultid="1659" />
                    <RANKING place="5" resultid="1772" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="7" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="7000" number="0" />
                <HEAT heatid="7001" number="1" />
                <HEAT heatid="7002" number="2" />
                <HEAT heatid="7003" number="3" />
                <HEAT heatid="7004" number="4" />
                <HEAT heatid="7005" number="5" />
                <HEAT heatid="7006" number="6" />
                <HEAT heatid="7007" number="7" />
                <HEAT heatid="7008" number="8" />
                <HEAT heatid="7009" number="9" />
                <HEAT heatid="7010" number="10" />
                <HEAT heatid="7011" number="11" />
                <HEAT heatid="7012" number="12" />
                <HEAT heatid="7013" number="13" />
                <HEAT heatid="7014" number="14" />
                <HEAT heatid="7015" number="15" />
                <HEAT heatid="7016" number="16" />
                <HEAT heatid="7017" number="17" />
                <HEAT heatid="7018" number="18" />
                <HEAT heatid="7019" number="19" />
                <HEAT heatid="7020" number="20" />
                <HEAT heatid="7021" number="21" />
                <HEAT heatid="7022" number="22" />
                <HEAT heatid="7023" number="23" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="12" resultid="303" />
                    <RANKING place="11" resultid="502" />
                    <RANKING place="2" resultid="538" />
                    <RANKING place="8" resultid="576" />
                    <RANKING place="1" resultid="580" />
                    <RANKING place="9" resultid="629" />
                    <RANKING place="3" resultid="641" />
                    <RANKING place="5" resultid="646" />
                    <RANKING place="4" resultid="790" />
                    <RANKING place="6" resultid="859" />
                    <RANKING place="7" resultid="1594" />
                    <RANKING place="13" resultid="1610" />
                    <RANKING place="10" resultid="1752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="7" resultid="356" />
                    <RANKING place="2" resultid="521" />
                    <RANKING place="5" resultid="687" />
                    <RANKING place="9" resultid="706" />
                    <RANKING place="12" resultid="759" />
                    <RANKING place="10" resultid="867" />
                    <RANKING place="3" resultid="955" />
                    <RANKING place="8" resultid="1291" />
                    <RANKING place="6" resultid="1299" />
                    <RANKING place="1" resultid="1302" />
                    <RANKING place="4" resultid="1502" />
                    <RANKING place="11" resultid="1518" />
                    <RANKING place="13" resultid="1903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="263" />
                    <RANKING place="14" resultid="446" />
                    <RANKING place="1" resultid="716" />
                    <RANKING place="3" resultid="748" />
                    <RANKING place="6" resultid="795" />
                    <RANKING place="4" resultid="812" />
                    <RANKING place="9" resultid="985" />
                    <RANKING place="12" resultid="1154" />
                    <RANKING place="16" resultid="1160" />
                    <RANKING place="7" resultid="1373" />
                    <RANKING place="15" resultid="1533" />
                    <RANKING place="10" resultid="1545" />
                    <RANKING place="5" resultid="1606" />
                    <RANKING place="13" resultid="1705" />
                    <RANKING place="11" resultid="1747" />
                    <RANKING place="8" resultid="1801" />
                    <RANKING place="17" resultid="1879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="7" resultid="275" />
                    <RANKING place="16" resultid="283" />
                    <RANKING place="17" resultid="470" />
                    <RANKING place="4" resultid="591" />
                    <RANKING place="13" resultid="722" />
                    <RANKING place="6" resultid="841" />
                    <RANKING place="12" resultid="1308" />
                    <RANKING place="8" resultid="1320" />
                    <RANKING place="1" resultid="1326" />
                    <RANKING place="3" resultid="1331" />
                    <RANKING place="14" resultid="1337" />
                    <RANKING place="2" resultid="1343" />
                    <RANKING place="11" resultid="1350" />
                    <RANKING place="9" resultid="1362" />
                    <RANKING place="5" resultid="1522" />
                    <RANKING place="15" resultid="1720" />
                    <RANKING place="10" resultid="1765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="10" resultid="50" />
                    <RANKING place="11" resultid="160" />
                    <RANKING place="8" resultid="271" />
                    <RANKING place="5" resultid="291" />
                    <RANKING place="2" resultid="414" />
                    <RANKING place="14" resultid="479" />
                    <RANKING place="7" resultid="526" />
                    <RANKING place="1" resultid="549" />
                    <RANKING place="6" resultid="564" />
                    <RANKING place="12" resultid="728" />
                    <RANKING place="9" resultid="1132" />
                    <RANKING place="17" resultid="1135" />
                    <RANKING place="15" resultid="1146" />
                    <RANKING place="16" resultid="1148" />
                    <RANKING place="18" resultid="1165" />
                    <RANKING place="19" resultid="1169" />
                    <RANKING place="4" resultid="1367" />
                    <RANKING place="22" resultid="1603" />
                    <RANKING place="13" resultid="1612" />
                    <RANKING place="3" resultid="1756" />
                    <RANKING place="20" resultid="1790" />
                    <RANKING place="21" resultid="1854" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="8" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="8000" number="0" />
                <HEAT heatid="8001" number="1" />
                <HEAT heatid="8002" number="2" />
                <HEAT heatid="8003" number="3" />
                <HEAT heatid="8004" number="4" />
                <HEAT heatid="8005" number="5" />
                <HEAT heatid="8006" number="6" />
                <HEAT heatid="8007" number="7" />
                <HEAT heatid="8008" number="8" />
                <HEAT heatid="8009" number="9" />
                <HEAT heatid="8010" number="10" />
                <HEAT heatid="8011" number="11" />
                <HEAT heatid="8012" number="12" />
                <HEAT heatid="8013" number="13" />
                <HEAT heatid="8014" number="14" />
                <HEAT heatid="8015" number="15" />
                <HEAT heatid="8016" number="16" />
                <HEAT heatid="8017" number="17" />
                <HEAT heatid="8018" number="18" />
                <HEAT heatid="8019" number="19" />
                <HEAT heatid="8020" number="20" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="672" />
                    <RANKING place="1" resultid="1379" />
                    <RANKING place="2" resultid="1897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="7" resultid="214" />
                    <RANKING place="9" resultid="237" />
                    <RANKING place="1" resultid="484" />
                    <RANKING place="3" resultid="488" />
                    <RANKING place="4" resultid="492" />
                    <RANKING place="6" resultid="650" />
                    <RANKING place="5" resultid="766" />
                    <RANKING place="8" resultid="908" />
                    <RANKING place="10" resultid="991" />
                    <RANKING place="2" resultid="1387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="431" />
                    <RANKING place="6" resultid="555" />
                    <RANKING place="8" resultid="623" />
                    <RANKING place="7" resultid="711" />
                    <RANKING place="17" resultid="886" />
                    <RANKING place="4" resultid="918" />
                    <RANKING place="19" resultid="1140" />
                    <RANKING place="13" resultid="1143" />
                    <RANKING place="2" resultid="1156" />
                    <RANKING place="9" resultid="1438" />
                    <RANKING place="5" resultid="1443" />
                    <RANKING place="3" resultid="1450" />
                    <RANKING place="10" resultid="1539" />
                    <RANKING place="14" resultid="1597" />
                    <RANKING place="12" resultid="1709" />
                    <RANKING place="20" resultid="1727" />
                    <RANKING place="17" resultid="1730" />
                    <RANKING place="11" resultid="1742" />
                    <RANKING place="16" resultid="1797" />
                    <RANKING place="15" resultid="1817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="14" resultid="362" />
                    <RANKING place="1" resultid="425" />
                    <RANKING place="2" resultid="698" />
                    <RANKING place="8" resultid="880" />
                    <RANKING place="5" resultid="1024" />
                    <RANKING place="16" resultid="1044" />
                    <RANKING place="6" resultid="1101" />
                    <RANKING place="13" resultid="1166" />
                    <RANKING place="12" resultid="1391" />
                    <RANKING place="7" resultid="1414" />
                    <RANKING place="9" resultid="1426" />
                    <RANKING place="10" resultid="1432" />
                    <RANKING place="3" resultid="1563" />
                    <RANKING place="4" resultid="1570" />
                    <RANKING place="11" resultid="1630" />
                    <RANKING place="15" resultid="1674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="5" resultid="340" />
                    <RANKING place="7" resultid="388" />
                    <RANKING place="2" resultid="532" />
                    <RANKING place="4" resultid="999" />
                    <RANKING place="9" resultid="1014" />
                    <RANKING place="3" resultid="1096" />
                    <RANKING place="8" resultid="1402" />
                    <RANKING place="10" resultid="1552" />
                    <RANKING place="1" resultid="1591" />
                    <RANKING place="11" resultid="1635" />
                    <RANKING place="6" resultid="1650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="4" resultid="33" />
                    <RANKING place="2" resultid="441" />
                    <RANKING place="6" resultid="543" />
                    <RANKING place="1" resultid="774" />
                    <RANKING place="5" resultid="830" />
                    <RANKING place="11" resultid="961" />
                    <RANKING place="9" resultid="1049" />
                    <RANKING place="8" resultid="1069" />
                    <RANKING place="3" resultid="1137" />
                    <RANKING place="10" resultid="1158" />
                    <RANKING place="7" resultid="1576" />
                    <RANKING place="12" resultid="1660" />
                    <RANKING place="13" resultid="1773" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="9" gender="F" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="9000" number="0" />
                <HEAT heatid="9001" number="1" />
                <HEAT heatid="9002" number="2" />
                <HEAT heatid="9003" number="3" />
                <HEAT heatid="9004" number="4" />
                <HEAT heatid="9005" number="5" />
                <HEAT heatid="9006" number="6" />
                <HEAT heatid="9007" number="7" />
                <HEAT heatid="9008" number="8" />
                <HEAT heatid="9009" number="9" />
                <HEAT heatid="9010" number="10" />
                <HEAT heatid="9011" number="11" />
                <HEAT heatid="9012" number="12" />
                <HEAT heatid="9013" number="13" />
                <HEAT heatid="9014" number="14" />
                <HEAT heatid="9015" number="15" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="539" />
                    <RANKING place="2" resultid="581" />
                    <RANKING place="1" resultid="642" />
                    <RANKING place="4" resultid="1595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="4" resultid="357" />
                    <RANKING place="9" resultid="518" />
                    <RANKING place="1" resultid="522" />
                    <RANKING place="5" resultid="619" />
                    <RANKING place="8" resultid="868" />
                    <RANKING place="7" resultid="956" />
                    <RANKING place="2" resultid="1295" />
                    <RANKING place="3" resultid="1303" />
                    <RANKING place="6" resultid="1503" />
                    <RANKING place="10" resultid="1519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="6" resultid="733" />
                    <RANKING place="3" resultid="796" />
                    <RANKING place="4" resultid="813" />
                    <RANKING place="1" resultid="937" />
                    <RANKING place="5" resultid="1374" />
                    <RANKING place="7" resultid="1491" />
                    <RANKING place="10" resultid="1534" />
                    <RANKING place="8" resultid="1546" />
                    <RANKING place="2" resultid="1607" />
                    <RANKING place="9" resultid="1706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="60" />
                    <RANKING place="9" resultid="241" />
                    <RANKING place="12" resultid="471" />
                    <RANKING place="4" resultid="592" />
                    <RANKING place="6" resultid="842" />
                    <RANKING place="2" resultid="1332" />
                    <RANKING place="10" resultid="1338" />
                    <RANKING place="1" resultid="1344" />
                    <RANKING place="5" resultid="1356" />
                    <RANKING place="7" resultid="1528" />
                    <RANKING place="11" resultid="1721" />
                    <RANKING place="8" resultid="1766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="9" resultid="36" />
                    <RANKING place="12" resultid="321" />
                    <RANKING place="10" resultid="480" />
                    <RANKING place="7" resultid="527" />
                    <RANKING place="5" resultid="565" />
                    <RANKING place="3" resultid="1055" />
                    <RANKING place="2" resultid="1368" />
                    <RANKING place="11" resultid="1601" />
                    <RANKING place="14" resultid="1604" />
                    <RANKING place="8" resultid="1613" />
                    <RANKING place="6" resultid="1692" />
                    <RANKING place="4" resultid="1757" />
                    <RANKING place="13" resultid="1791" />
                    <RANKING place="15" resultid="1855" />
                    <RANKING place="1" resultid="1866" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="10" number="10" gender="M" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="10000" number="0" />
                <HEAT heatid="10001" number="1" />
                <HEAT heatid="10002" number="2" />
                <HEAT heatid="10003" number="3" />
                <HEAT heatid="10004" number="4" />
                <HEAT heatid="10005" number="5" />
                <HEAT heatid="10006" number="6" />
                <HEAT heatid="10007" number="7" />
                <HEAT heatid="10008" number="8" />
                <HEAT heatid="10009" number="9" />
                <HEAT heatid="10010" number="10" />
                <HEAT heatid="10011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="2" resultid="673" />
                    <RANKING place="1" resultid="1898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="6" resultid="215" />
                    <RANKING place="1" resultid="651" />
                    <RANKING place="2" resultid="767" />
                    <RANKING place="3" resultid="909" />
                    <RANKING place="5" resultid="992" />
                    <RANKING place="4" resultid="1654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="249" />
                    <RANKING place="6" resultid="299" />
                    <RANKING place="7" resultid="624" />
                    <RANKING place="8" resultid="712" />
                    <RANKING place="5" resultid="919" />
                    <RANKING place="3" resultid="1444" />
                    <RANKING place="1" resultid="1456" />
                    <RANKING place="4" resultid="1540" />
                    <RANKING place="10" resultid="1598" />
                    <RANKING place="9" resultid="1710" />
                    <RANKING place="11" resultid="1731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="9" />
                    <RANKING place="4" resultid="15" />
                    <RANKING place="3" resultid="21" />
                    <RANKING place="7" resultid="363" />
                    <RANKING place="2" resultid="699" />
                    <RANKING place="8" resultid="1045" />
                    <RANKING place="5" resultid="1102" />
                    <RANKING place="6" resultid="1564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="341" />
                    <RANKING place="2" resultid="1015" />
                    <RANKING place="1" resultid="1592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="442" />
                    <RANKING place="6" resultid="544" />
                    <RANKING place="1" resultid="775" />
                    <RANKING place="4" resultid="831" />
                    <RANKING place="7" resultid="1050" />
                    <RANKING place="5" resultid="1070" />
                    <RANKING place="3" resultid="1138" />
                    <RANKING place="8" resultid="1661" />
                    <RANKING place="9" resultid="1774" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="11" gender="X" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="11001" number="1" />
                <HEAT heatid="11002" number="2" />
                <HEAT heatid="11003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="13" agemin="8" name="Jahrgänge 2010 bis 2015">
                  <RANKINGS>
                    <RANKING place="2" resultid="260" />
                    <RANKING place="10" resultid="309" />
                    <RANKING place="1" resultid="495" />
                    <RANKING place="3" resultid="787" />
                    <RANKING place="5" resultid="1466" />
                    <RANKING place="7" resultid="1468" />
                    <RANKING place="4" resultid="1488" />
                    <RANKING place="6" resultid="1618" />
                    <RANKING place="9" resultid="1624" />
                    <RANKING place="8" resultid="1958" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2023-12-09" daytime="14:00">
          <EVENTS>
            <EVENT eventid="13" number="12" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="13000" number="0" />
                <HEAT heatid="13001" number="1" />
                <HEAT heatid="13002" number="2" />
                <HEAT heatid="13003" number="3" />
                <HEAT heatid="13004" number="4" />
                <HEAT heatid="13005" number="5" />
                <HEAT heatid="13006" number="6" />
                <HEAT heatid="13007" number="7" />
                <HEAT heatid="13008" number="8" />
                <HEAT heatid="13009" number="9" />
                <HEAT heatid="13010" number="10" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="1" resultid="582" />
                    <RANKING place="2" resultid="643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="523" />
                    <RANKING place="5" resultid="869" />
                    <RANKING place="4" resultid="957" />
                    <RANKING place="3" resultid="1304" />
                    <RANKING place="2" resultid="1504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="717" />
                    <RANKING place="2" resultid="749" />
                    <RANKING place="3" resultid="814" />
                    <RANKING place="4" resultid="1492" />
                    <RANKING place="6" resultid="1535" />
                    <RANKING place="5" resultid="1547" />
                    <RANKING place="7" resultid="1748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="9" resultid="242" />
                    <RANKING place="13" resultid="284" />
                    <RANKING place="1" resultid="593" />
                    <RANKING place="11" resultid="723" />
                    <RANKING place="2" resultid="843" />
                    <RANKING place="3" resultid="1327" />
                    <RANKING place="4" resultid="1333" />
                    <RANKING place="12" resultid="1339" />
                    <RANKING place="5" resultid="1345" />
                    <RANKING place="10" resultid="1351" />
                    <RANKING place="7" resultid="1357" />
                    <RANKING place="6" resultid="1523" />
                    <RANKING place="8" resultid="1529" />
                    <RANKING place="14" resultid="1722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="5" resultid="37" />
                    <RANKING place="2" resultid="528" />
                    <RANKING place="1" resultid="550" />
                    <RANKING place="4" resultid="1693" />
                    <RANKING place="3" resultid="1758" />
                    <RANKING place="6" resultid="1792" />
                    <RANKING place="7" resultid="1856" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="14" number="13" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="14000" number="0" />
                <HEAT heatid="14001" number="1" />
                <HEAT heatid="14002" number="2" />
                <HEAT heatid="14003" number="3" />
                <HEAT heatid="14004" number="4" />
                <HEAT heatid="14005" number="5" />
                <HEAT heatid="14006" number="6" />
                <HEAT heatid="14007" number="7" />
                <HEAT heatid="14008" number="8" />
                <HEAT heatid="14009" number="9" />
                <HEAT heatid="14010" number="10" />
                <HEAT heatid="14011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="1" resultid="1380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="485" />
                    <RANKING place="4" resultid="768" />
                    <RANKING place="2" resultid="1388" />
                    <RANKING place="3" resultid="1655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="6" resultid="250" />
                    <RANKING place="7" resultid="300" />
                    <RANKING place="2" resultid="432" />
                    <RANKING place="9" resultid="556" />
                    <RANKING place="8" resultid="713" />
                    <RANKING place="1" resultid="1445" />
                    <RANKING place="3" resultid="1451" />
                    <RANKING place="4" resultid="1457" />
                    <RANKING place="5" resultid="1541" />
                    <RANKING place="11" resultid="1711" />
                    <RANKING place="10" resultid="1732" />
                    <RANKING place="12" resultid="1743" />
                    <RANKING place="13" resultid="1818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="10" />
                    <RANKING place="2" resultid="307" />
                    <RANKING place="3" resultid="700" />
                    <RANKING place="7" resultid="881" />
                    <RANKING place="4" resultid="1025" />
                    <RANKING place="6" resultid="1565" />
                    <RANKING place="5" resultid="1571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="342" />
                    <RANKING place="5" resultid="390" />
                    <RANKING place="1" resultid="533" />
                    <RANKING place="2" resultid="1000" />
                    <RANKING place="3" resultid="1097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="443" />
                    <RANKING place="1" resultid="776" />
                    <RANKING place="3" resultid="1151" />
                    <RANKING place="4" resultid="1577" />
                    <RANKING place="5" resultid="1662" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="15" number="14" gender="F" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="15000" number="0" />
                <HEAT heatid="15001" number="1" />
                <HEAT heatid="15002" number="2" />
                <HEAT heatid="15003" number="3" />
                <HEAT heatid="15004" number="4" />
                <HEAT heatid="15005" number="5" />
                <HEAT heatid="15006" number="6" />
                <HEAT heatid="15007" number="7" />
                <HEAT heatid="15008" number="8" />
                <HEAT heatid="15009" number="9" />
                <HEAT heatid="15010" number="10" />
                <HEAT heatid="15011" number="11" />
                <HEAT heatid="15012" number="12" />
                <HEAT heatid="15013" number="13" />
                <HEAT heatid="15014" number="14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="5" resultid="503" />
                    <RANKING place="2" resultid="540" />
                    <RANKING place="6" resultid="647" />
                    <RANKING place="1" resultid="791" />
                    <RANKING place="3" resultid="802" />
                    <RANKING place="4" resultid="1514" />
                    <RANKING place="7" resultid="1753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="4" resultid="358" />
                    <RANKING place="6" resultid="587" />
                    <RANKING place="5" resultid="688" />
                    <RANKING place="2" resultid="958" />
                    <RANKING place="3" resultid="1292" />
                    <RANKING place="1" resultid="1296" />
                    <RANKING place="7" resultid="1904" />
                    <RANKING place="8" resultid="1928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="264" />
                    <RANKING place="8" resultid="448" />
                    <RANKING place="1" resultid="718" />
                    <RANKING place="3" resultid="797" />
                    <RANKING place="4" resultid="815" />
                    <RANKING place="6" resultid="987" />
                    <RANKING place="5" resultid="1375" />
                    <RANKING place="10" resultid="1536" />
                    <RANKING place="9" resultid="1749" />
                    <RANKING place="7" resultid="1802" />
                    <RANKING place="11" resultid="1881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="7" resultid="243" />
                    <RANKING place="3" resultid="276" />
                    <RANKING place="12" resultid="285" />
                    <RANKING place="8" resultid="724" />
                    <RANKING place="6" resultid="1309" />
                    <RANKING place="4" resultid="1321" />
                    <RANKING place="2" resultid="1328" />
                    <RANKING place="1" resultid="1334" />
                    <RANKING place="9" resultid="1340" />
                    <RANKING place="10" resultid="1363" />
                    <RANKING place="5" resultid="1524" />
                    <RANKING place="11" resultid="1767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="7" resultid="161" />
                    <RANKING place="9" resultid="272" />
                    <RANKING place="4" resultid="292" />
                    <RANKING place="2" resultid="415" />
                    <RANKING place="11" resultid="481" />
                    <RANKING place="1" resultid="551" />
                    <RANKING place="3" resultid="566" />
                    <RANKING place="8" resultid="729" />
                    <RANKING place="6" resultid="1369" />
                    <RANKING place="10" resultid="1694" />
                    <RANKING place="12" resultid="1793" />
                    <RANKING place="5" resultid="1867" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="16" number="15" gender="M" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="16000" number="0" />
                <HEAT heatid="16001" number="1" />
                <HEAT heatid="16002" number="2" />
                <HEAT heatid="16003" number="3" />
                <HEAT heatid="16004" number="4" />
                <HEAT heatid="16005" number="5" />
                <HEAT heatid="16006" number="6" />
                <HEAT heatid="16007" number="7" />
                <HEAT heatid="16008" number="8" />
                <HEAT heatid="16009" number="9" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="1" resultid="674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="238" />
                    <RANKING place="1" resultid="652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="6" resultid="557" />
                    <RANKING place="2" resultid="625" />
                    <RANKING place="5" resultid="921" />
                    <RANKING place="4" resultid="1439" />
                    <RANKING place="3" resultid="1446" />
                    <RANKING place="1" resultid="1452" />
                    <RANKING place="7" resultid="1744" />
                    <RANKING place="8" resultid="1819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="16" />
                    <RANKING place="4" resultid="426" />
                    <RANKING place="1" resultid="701" />
                    <RANKING place="2" resultid="1026" />
                    <RANKING place="6" resultid="1103" />
                    <RANKING place="5" resultid="1415" />
                    <RANKING place="9" resultid="1427" />
                    <RANKING place="8" resultid="1433" />
                    <RANKING place="7" resultid="1566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="534" />
                    <RANKING place="2" resultid="1016" />
                    <RANKING place="3" resultid="1403" />
                    <RANKING place="5" resultid="1553" />
                    <RANKING place="4" resultid="1651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="4" resultid="545" />
                    <RANKING place="2" resultid="832" />
                    <RANKING place="5" resultid="963" />
                    <RANKING place="1" resultid="1071" />
                    <RANKING place="3" resultid="1578" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="17" number="16" gender="F" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="17000" number="0" />
                <HEAT heatid="17001" number="1" />
                <HEAT heatid="17002" number="2" />
                <HEAT heatid="17003" number="3" />
                <HEAT heatid="17004" number="4" />
                <HEAT heatid="17005" number="5" />
                <HEAT heatid="17006" number="6" />
                <HEAT heatid="17007" number="7" />
                <HEAT heatid="17008" number="8" />
                <HEAT heatid="17009" number="9" />
                <HEAT heatid="17010" number="10" />
                <HEAT heatid="17011" number="11" />
                <HEAT heatid="17012" number="12" />
                <HEAT heatid="17013" number="13" />
                <HEAT heatid="17014" number="14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="9" resultid="304" />
                    <RANKING place="10" resultid="504" />
                    <RANKING place="6" resultid="577" />
                    <RANKING place="2" resultid="583" />
                    <RANKING place="7" resultid="630" />
                    <RANKING place="1" resultid="792" />
                    <RANKING place="5" resultid="803" />
                    <RANKING place="8" resultid="860" />
                    <RANKING place="4" resultid="1515" />
                    <RANKING place="3" resultid="1754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="6" resultid="519" />
                    <RANKING place="2" resultid="588" />
                    <RANKING place="5" resultid="620" />
                    <RANKING place="1" resultid="689" />
                    <RANKING place="4" resultid="708" />
                    <RANKING place="8" resultid="760" />
                    <RANKING place="3" resultid="870" />
                    <RANKING place="7" resultid="1905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="694" />
                    <RANKING place="7" resultid="734" />
                    <RANKING place="1" resultid="939" />
                    <RANKING place="9" resultid="988" />
                    <RANKING place="11" resultid="1155" />
                    <RANKING place="12" resultid="1161" />
                    <RANKING place="5" resultid="1376" />
                    <RANKING place="8" resultid="1493" />
                    <RANKING place="3" resultid="1548" />
                    <RANKING place="4" resultid="1707" />
                    <RANKING place="6" resultid="1803" />
                    <RANKING place="10" resultid="1882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="61" />
                    <RANKING place="10" resultid="772" />
                    <RANKING place="6" resultid="1310" />
                    <RANKING place="8" resultid="1322" />
                    <RANKING place="3" resultid="1352" />
                    <RANKING place="1" resultid="1358" />
                    <RANKING place="5" resultid="1364" />
                    <RANKING place="4" resultid="1530" />
                    <RANKING place="9" resultid="1723" />
                    <RANKING place="7" resultid="1768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="5" resultid="567" />
                    <RANKING place="8" resultid="730" />
                    <RANKING place="1" resultid="1056" />
                    <RANKING place="2" resultid="1133" />
                    <RANKING place="9" resultid="1136" />
                    <RANKING place="6" resultid="1370" />
                    <RANKING place="3" resultid="1695" />
                    <RANKING place="7" resultid="1759" />
                    <RANKING place="10" resultid="1857" />
                    <RANKING place="4" resultid="1868" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18" number="17" gender="M" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="18000" number="0" />
                <HEAT heatid="18001" number="1" />
                <HEAT heatid="18002" number="2" />
                <HEAT heatid="18003" number="3" />
                <HEAT heatid="18004" number="4" />
                <HEAT heatid="18005" number="5" />
                <HEAT heatid="18006" number="6" />
                <HEAT heatid="18007" number="7" />
                <HEAT heatid="18008" number="8" />
                <HEAT heatid="18009" number="9" />
                <HEAT heatid="18010" number="10" />
                <HEAT heatid="18011" number="11" />
                <HEAT heatid="18012" number="12" />
                <HEAT heatid="18013" number="13" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="2" resultid="675" />
                    <RANKING place="1" resultid="1899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="653" />
                    <RANKING place="2" resultid="769" />
                    <RANKING place="3" resultid="910" />
                    <RANKING place="4" resultid="1656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="251" />
                    <RANKING place="2" resultid="714" />
                    <RANKING place="7" resultid="887" />
                    <RANKING place="5" resultid="1144" />
                    <RANKING place="4" resultid="1440" />
                    <RANKING place="6" resultid="1542" />
                    <RANKING place="3" resultid="1712" />
                    <RANKING place="8" resultid="1728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="17" />
                    <RANKING place="1" resultid="22" />
                    <RANKING place="12" resultid="364" />
                    <RANKING place="3" resultid="882" />
                    <RANKING place="11" resultid="1046" />
                    <RANKING place="5" resultid="1167" />
                    <RANKING place="6" resultid="1416" />
                    <RANKING place="9" resultid="1428" />
                    <RANKING place="8" resultid="1434" />
                    <RANKING place="4" resultid="1572" />
                    <RANKING place="10" resultid="1632" />
                    <RANKING place="7" resultid="1675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="5" resultid="391" />
                    <RANKING place="2" resultid="1001" />
                    <RANKING place="1" resultid="1098" />
                    <RANKING place="4" resultid="1404" />
                    <RANKING place="6" resultid="1554" />
                    <RANKING place="3" resultid="1636" />
                    <RANKING place="7" resultid="1652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="7" resultid="546" />
                    <RANKING place="1" resultid="777" />
                    <RANKING place="3" resultid="833" />
                    <RANKING place="6" resultid="1051" />
                    <RANKING place="8" resultid="1072" />
                    <RANKING place="2" resultid="1152" />
                    <RANKING place="4" resultid="1579" />
                    <RANKING place="5" resultid="1663" />
                    <RANKING place="9" resultid="1775" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="19" number="18" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="19000" number="0" />
                <HEAT heatid="19001" number="1" />
                <HEAT heatid="19002" number="2" />
                <HEAT heatid="19003" number="3" />
                <HEAT heatid="19004" number="4" />
                <HEAT heatid="19005" number="5" />
                <HEAT heatid="19006" number="6" />
                <HEAT heatid="19007" number="7" />
                <HEAT heatid="19008" number="8" />
                <HEAT heatid="19009" number="9" />
                <HEAT heatid="19010" number="10" />
                <HEAT heatid="19011" number="11" />
                <HEAT heatid="19012" number="12" />
                <HEAT heatid="19013" number="13" />
                <HEAT heatid="19014" number="14" />
                <HEAT heatid="19015" number="15" />
                <HEAT heatid="19016" number="16" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="541" />
                    <RANKING place="8" resultid="578" />
                    <RANKING place="1" resultid="584" />
                    <RANKING place="4" resultid="631" />
                    <RANKING place="6" resultid="648" />
                    <RANKING place="2" resultid="793" />
                    <RANKING place="7" resultid="861" />
                    <RANKING place="5" resultid="1516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="8" resultid="359" />
                    <RANKING place="3" resultid="524" />
                    <RANKING place="12" resultid="589" />
                    <RANKING place="10" resultid="621" />
                    <RANKING place="4" resultid="690" />
                    <RANKING place="9" resultid="871" />
                    <RANKING place="11" resultid="959" />
                    <RANKING place="7" resultid="1293" />
                    <RANKING place="1" resultid="1297" />
                    <RANKING place="6" resultid="1301" />
                    <RANKING place="2" resultid="1305" />
                    <RANKING place="5" resultid="1506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="265" />
                    <RANKING place="12" resultid="449" />
                    <RANKING place="8" resultid="695" />
                    <RANKING place="1" resultid="719" />
                    <RANKING place="9" resultid="735" />
                    <RANKING place="3" resultid="750" />
                    <RANKING place="4" resultid="798" />
                    <RANKING place="5" resultid="816" />
                    <RANKING place="7" resultid="989" />
                    <RANKING place="6" resultid="1377" />
                    <RANKING place="11" resultid="1494" />
                    <RANKING place="14" resultid="1537" />
                    <RANKING place="10" resultid="1549" />
                    <RANKING place="13" resultid="1804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="62" />
                    <RANKING place="16" resultid="472" />
                    <RANKING place="2" resultid="594" />
                    <RANKING place="15" resultid="725" />
                    <RANKING place="6" resultid="844" />
                    <RANKING place="12" resultid="1311" />
                    <RANKING place="5" resultid="1323" />
                    <RANKING place="7" resultid="1329" />
                    <RANKING place="3" resultid="1335" />
                    <RANKING place="14" resultid="1341" />
                    <RANKING place="1" resultid="1346" />
                    <RANKING place="10" resultid="1353" />
                    <RANKING place="9" resultid="1365" />
                    <RANKING place="11" resultid="1525" />
                    <RANKING place="8" resultid="1531" />
                    <RANKING place="13" resultid="1769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="10" resultid="322" />
                    <RANKING place="2" resultid="416" />
                    <RANKING place="7" resultid="482" />
                    <RANKING place="1" resultid="552" />
                    <RANKING place="5" resultid="568" />
                    <RANKING place="3" resultid="1057" />
                    <RANKING place="8" resultid="1149" />
                    <RANKING place="6" resultid="1371" />
                    <RANKING place="4" resultid="1760" />
                    <RANKING place="9" resultid="1794" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="20" number="19" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="20000" number="0" />
                <HEAT heatid="20001" number="1" />
                <HEAT heatid="20002" number="2" />
                <HEAT heatid="20003" number="3" />
                <HEAT heatid="20004" number="4" />
                <HEAT heatid="20005" number="5" />
                <HEAT heatid="20006" number="6" />
                <HEAT heatid="20007" number="7" />
                <HEAT heatid="20008" number="8" />
                <HEAT heatid="20009" number="9" />
                <HEAT heatid="20010" number="10" />
                <HEAT heatid="20011" number="11" />
                <HEAT heatid="20012" number="12" />
                <HEAT heatid="20013" number="13" />
                <HEAT heatid="20014" number="14" />
                <HEAT heatid="20015" number="15" />
                <HEAT heatid="20016" number="16" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="676" />
                    <RANKING place="1" resultid="1381" />
                    <RANKING place="2" resultid="1900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="6" resultid="217" />
                    <RANKING place="8" resultid="239" />
                    <RANKING place="1" resultid="486" />
                    <RANKING place="3" resultid="494" />
                    <RANKING place="4" resultid="654" />
                    <RANKING place="5" resultid="911" />
                    <RANKING place="9" resultid="993" />
                    <RANKING place="2" resultid="1389" />
                    <RANKING place="7" resultid="1657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="8" resultid="301" />
                    <RANKING place="1" resultid="433" />
                    <RANKING place="9" resultid="558" />
                    <RANKING place="5" resultid="626" />
                    <RANKING place="15" resultid="888" />
                    <RANKING place="6" resultid="922" />
                    <RANKING place="3" resultid="1157" />
                    <RANKING place="7" resultid="1441" />
                    <RANKING place="4" resultid="1447" />
                    <RANKING place="2" resultid="1453" />
                    <RANKING place="10" resultid="1543" />
                    <RANKING place="12" resultid="1733" />
                    <RANKING place="11" resultid="1745" />
                    <RANKING place="14" resultid="1799" />
                    <RANKING place="13" resultid="1820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="308" />
                    <RANKING place="13" resultid="365" />
                    <RANKING place="2" resultid="427" />
                    <RANKING place="3" resultid="702" />
                    <RANKING place="9" resultid="883" />
                    <RANKING place="7" resultid="1027" />
                    <RANKING place="14" resultid="1047" />
                    <RANKING place="8" resultid="1104" />
                    <RANKING place="12" resultid="1393" />
                    <RANKING place="6" resultid="1417" />
                    <RANKING place="11" resultid="1429" />
                    <RANKING place="10" resultid="1435" />
                    <RANKING place="4" resultid="1567" />
                    <RANKING place="5" resultid="1573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="343" />
                    <RANKING place="1" resultid="535" />
                    <RANKING place="3" resultid="1002" />
                    <RANKING place="4" resultid="1017" />
                    <RANKING place="2" resultid="1099" />
                    <RANKING place="5" resultid="1405" />
                    <RANKING place="8" resultid="1555" />
                    <RANKING place="9" resultid="1637" />
                    <RANKING place="7" resultid="1653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="444" />
                    <RANKING place="1" resultid="778" />
                    <RANKING place="4" resultid="834" />
                    <RANKING place="6" resultid="964" />
                    <RANKING place="5" resultid="1052" />
                    <RANKING place="3" resultid="1139" />
                    <RANKING place="7" resultid="1664" />
                    <RANKING place="8" resultid="1776" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="21" number="20" gender="F" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="21001" number="1" />
                <HEAT heatid="21002" number="2" />
                <HEAT heatid="21003" number="3" />
                <HEAT heatid="21004" number="4" />
                <HEAT heatid="21005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="720" />
                    <RANKING place="4" resultid="751" />
                    <RANKING place="3" resultid="799" />
                    <RANKING place="1" resultid="940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="277" />
                    <RANKING place="3" resultid="595" />
                    <RANKING place="4" resultid="845" />
                    <RANKING place="1" resultid="1347" />
                    <RANKING place="5" resultid="1359" />
                    <RANKING place="6" resultid="1724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="51" />
                    <RANKING place="5" resultid="162" />
                    <RANKING place="4" resultid="273" />
                    <RANKING place="3" resultid="293" />
                    <RANKING place="1" resultid="553" />
                    <RANKING place="2" resultid="1869" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22" number="21" gender="M" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="22000" number="0" />
                <HEAT heatid="22001" number="1" />
                <HEAT heatid="22002" number="2" />
                <HEAT heatid="22003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="627" />
                    <RANKING place="2" resultid="1713" />
                    <RANKING place="3" resultid="1734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="12" agemin="12" name="Jahrgang 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="34" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23" number="22" gender="X" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="23001" number="1" />
                <HEAT heatid="23002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="13" agemin="8" name="Jahrgänge 2010 bis 2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="261" />
                    <RANKING place="5" resultid="310" />
                    <RANKING place="1" resultid="496" />
                    <RANKING place="2" resultid="788" />
                    <RANKING place="6" resultid="1467" />
                    <RANKING place="8" resultid="1469" />
                    <RANKING place="4" resultid="1619" />
                    <RANKING place="7" resultid="1625" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="3" date="2023-12-10" daytime="08:45" officialmeeting="08:15" warmupfrom="07:30">
          <EVENTS>
            <EVENT eventid="25" number="23" gender="F" round="PRE">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="25000" number="0" />
                <HEAT heatid="25001" number="1" />
                <HEAT heatid="25002" number="2" />
                <HEAT heatid="25003" number="3" />
                <HEAT heatid="25004" number="4" />
                <HEAT heatid="25005" number="5" />
                <HEAT heatid="25006" number="6" />
                <HEAT heatid="25007" number="7" />
                <HEAT heatid="25008" number="8" />
                <HEAT heatid="25009" number="9" />
                <HEAT heatid="25010" number="10" />
                <HEAT heatid="25011" number="11" />
                <HEAT heatid="25012" number="12" />
                <HEAT heatid="25013" number="13" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="3" resultid="367" />
                    <RANKING place="5" resultid="569" />
                    <RANKING place="2" resultid="923" />
                    <RANKING place="1" resultid="1008" />
                    <RANKING place="4" resultid="1665" />
                    <RANKING place="6" resultid="1735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="5" resultid="464" />
                    <RANKING place="6" resultid="505" />
                    <RANKING place="2" resultid="602" />
                    <RANKING place="3" resultid="741" />
                    <RANKING place="1" resultid="872" />
                    <RANKING place="4" resultid="1028" />
                    <RANKING place="6" resultid="1038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="17" resultid="163" />
                    <RANKING place="11" resultid="184" />
                    <RANKING place="2" resultid="266" />
                    <RANKING place="12" resultid="596" />
                    <RANKING place="5" resultid="667" />
                    <RANKING place="8" resultid="779" />
                    <RANKING place="14" resultid="835" />
                    <RANKING place="16" resultid="941" />
                    <RANKING place="18" resultid="1105" />
                    <RANKING place="19" resultid="1126" />
                    <RANKING place="6" resultid="1179" />
                    <RANKING place="15" resultid="1183" />
                    <RANKING place="9" resultid="1189" />
                    <RANKING place="1" resultid="1203" />
                    <RANKING place="7" resultid="1223" />
                    <RANKING place="4" resultid="1235" />
                    <RANKING place="2" resultid="1240" />
                    <RANKING place="22" resultid="1685" />
                    <RANKING place="20" resultid="1714" />
                    <RANKING place="13" resultid="1847" />
                    <RANKING place="21" resultid="1858" />
                    <RANKING place="10" resultid="1872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="2" resultid="52" />
                    <RANKING place="1" resultid="419" />
                    <RANKING place="3" resultid="752" />
                    <RANKING place="4" resultid="912" />
                    <RANKING place="5" resultid="1906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="148" />
                    <RANKING place="5" resultid="900" />
                    <RANKING place="7" resultid="965" />
                    <RANKING place="6" resultid="1584" />
                    <RANKING place="4" resultid="1698" />
                    <RANKING place="1" resultid="1807" />
                    <RANKING place="3" resultid="1840" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26" number="24" gender="M" round="PRE">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="26000" number="0" />
                <HEAT heatid="26001" number="1" />
                <HEAT heatid="26002" number="2" />
                <HEAT heatid="26003" number="3" />
                <HEAT heatid="26004" number="4" />
                <HEAT heatid="26005" number="5" />
                <HEAT heatid="26006" number="6" />
                <HEAT heatid="26007" number="7" />
                <HEAT heatid="26008" number="8" />
                <HEAT heatid="26009" number="9" />
                <HEAT heatid="26010" number="10" />
                <HEAT heatid="26011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="8" resultid="38" />
                    <RANKING place="4" resultid="374" />
                    <RANKING place="9" resultid="736" />
                    <RANKING place="5" resultid="889" />
                    <RANKING place="2" resultid="948" />
                    <RANKING place="7" resultid="1274" />
                    <RANKING place="1" resultid="1638" />
                    <RANKING place="6" resultid="1777" />
                    <RANKING place="10" resultid="1888" />
                    <RANKING place="3" resultid="1940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="10" resultid="153" />
                    <RANKING place="7" resultid="218" />
                    <RANKING place="3" resultid="278" />
                    <RANKING place="12" resultid="344" />
                    <RANKING place="8" resultid="398" />
                    <RANKING place="4" resultid="608" />
                    <RANKING place="6" resultid="677" />
                    <RANKING place="11" resultid="1078" />
                    <RANKING place="5" resultid="1254" />
                    <RANKING place="1" resultid="1263" />
                    <RANKING place="9" resultid="1676" />
                    <RANKING place="2" resultid="1834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="9" resultid="393" />
                    <RANKING place="3" resultid="632" />
                    <RANKING place="1" resultid="851" />
                    <RANKING place="7" resultid="1058" />
                    <RANKING place="2" resultid="1268" />
                    <RANKING place="4" resultid="1285" />
                    <RANKING place="8" resultid="1478" />
                    <RANKING place="6" resultid="1481" />
                    <RANKING place="5" resultid="1915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="655" />
                    <RANKING place="8" resultid="894" />
                    <RANKING place="3" resultid="930" />
                    <RANKING place="7" resultid="972" />
                    <RANKING place="6" resultid="1119" />
                    <RANKING place="2" resultid="1170" />
                    <RANKING place="5" resultid="1259" />
                    <RANKING place="1" resultid="1811" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="27" number="25" gender="F" round="PRE">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="27000" number="0" />
                <HEAT heatid="27001" number="1" />
                <HEAT heatid="27002" number="2" />
                <HEAT heatid="27003" number="3" />
                <HEAT heatid="27004" number="4" />
                <HEAT heatid="27005" number="5" />
                <HEAT heatid="27006" number="6" />
                <HEAT heatid="27007" number="7" />
                <HEAT heatid="27008" number="8" />
                <HEAT heatid="27009" number="9" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="29" />
                    <RANKING place="1" resultid="334" />
                    <RANKING place="4" resultid="570" />
                    <RANKING place="3" resultid="1018" />
                    <RANKING place="6" resultid="1033" />
                    <RANKING place="5" resultid="1073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="5" resultid="465" />
                    <RANKING place="8" resultid="506" />
                    <RANKING place="3" resultid="742" />
                    <RANKING place="2" resultid="873" />
                    <RANKING place="4" resultid="1085" />
                    <RANKING place="7" resultid="1121" />
                    <RANKING place="6" resultid="1557" />
                    <RANKING place="1" resultid="1929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="5" resultid="203" />
                    <RANKING place="3" resultid="256" />
                    <RANKING place="2" resultid="668" />
                    <RANKING place="6" resultid="836" />
                    <RANKING place="8" resultid="942" />
                    <RANKING place="1" resultid="1180" />
                    <RANKING place="4" resultid="1184" />
                    <RANKING place="7" resultid="1873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="3" resultid="53" />
                    <RANKING place="2" resultid="143" />
                    <RANKING place="1" resultid="1228" />
                    <RANKING place="4" resultid="1907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="169" />
                    <RANKING place="2" resultid="823" />
                    <RANKING place="4" resultid="862" />
                    <RANKING place="3" resultid="1585" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="28" number="26" gender="M" round="PRE">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="28000" number="0" />
                <HEAT heatid="28001" number="1" />
                <HEAT heatid="28002" number="2" />
                <HEAT heatid="28003" number="3" />
                <HEAT heatid="28004" number="4" />
                <HEAT heatid="28005" number="5" />
                <HEAT heatid="28006" number="6" />
                <HEAT heatid="28007" number="7" />
                <HEAT heatid="28008" number="8" />
                <HEAT heatid="28009" number="9" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="2" resultid="69" />
                    <RANKING place="1" resultid="375" />
                    <RANKING place="4" resultid="473" />
                    <RANKING place="6" resultid="737" />
                    <RANKING place="5" resultid="1275" />
                    <RANKING place="3" resultid="1639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="10" resultid="198" />
                    <RANKING place="9" resultid="219" />
                    <RANKING place="5" resultid="223" />
                    <RANKING place="11" resultid="399" />
                    <RANKING place="16" resultid="455" />
                    <RANKING place="8" resultid="609" />
                    <RANKING place="1" resultid="678" />
                    <RANKING place="13" resultid="1003" />
                    <RANKING place="7" resultid="1063" />
                    <RANKING place="2" resultid="1264" />
                    <RANKING place="12" resultid="1495" />
                    <RANKING place="6" resultid="1507" />
                    <RANKING place="4" resultid="1677" />
                    <RANKING place="13" resultid="1783" />
                    <RANKING place="3" resultid="1835" />
                    <RANKING place="15" resultid="1951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="5" resultid="394" />
                    <RANKING place="6" resultid="407" />
                    <RANKING place="2" resultid="852" />
                    <RANKING place="3" resultid="1090" />
                    <RANKING place="1" resultid="1269" />
                    <RANKING place="7" resultid="1821" />
                    <RANKING place="8" resultid="1827" />
                    <RANKING place="4" resultid="1916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="380" />
                    <RANKING place="5" resultid="895" />
                    <RANKING place="3" resultid="931" />
                    <RANKING place="2" resultid="1202" />
                    <RANKING place="1" resultid="1812" />
                    <RANKING place="6" resultid="1921" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="29" number="27" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="29000" number="0" />
                <HEAT heatid="29001" number="1" />
                <HEAT heatid="29002" number="2" />
                <HEAT heatid="29003" number="3" />
                <HEAT heatid="29004" number="4" />
                <HEAT heatid="29005" number="5" />
                <HEAT heatid="29006" number="6" />
                <HEAT heatid="29007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="5" resultid="41" />
                    <RANKING place="2" resultid="924" />
                    <RANKING place="1" resultid="1009" />
                    <RANKING place="4" resultid="1246" />
                    <RANKING place="3" resultid="1666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="1" resultid="603" />
                    <RANKING place="2" resultid="1930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="1" resultid="193" />
                    <RANKING place="2" resultid="267" />
                    <RANKING place="4" resultid="780" />
                    <RANKING place="6" resultid="1106" />
                    <RANKING place="5" resultid="1127" />
                    <RANKING place="3" resultid="1198" />
                    <RANKING place="7" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="3" resultid="189" />
                    <RANKING place="1" resultid="753" />
                    <RANKING place="2" resultid="1114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="149" />
                    <RANKING place="4" resultid="824" />
                    <RANKING place="3" resultid="901" />
                    <RANKING place="5" resultid="966" />
                    <RANKING place="2" resultid="1841" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="30" number="28" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="30001" number="1" />
                <HEAT heatid="30002" number="2" />
                <HEAT heatid="30003" number="3" />
                <HEAT heatid="30004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="2" resultid="228" />
                    <RANKING place="3" resultid="949" />
                    <RANKING place="1" resultid="1640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="179" />
                    <RANKING place="2" resultid="610" />
                    <RANKING place="5" resultid="1064" />
                    <RANKING place="4" resultid="1255" />
                    <RANKING place="1" resultid="1279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="1" resultid="633" />
                    <RANKING place="2" resultid="1828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="85" />
                    <RANKING place="3" resultid="381" />
                    <RANKING place="4" resultid="656" />
                    <RANKING place="2" resultid="896" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="31" number="29" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="31000" number="0" />
                <HEAT heatid="31001" number="1" />
                <HEAT heatid="31002" number="2" />
                <HEAT heatid="31003" number="3" />
                <HEAT heatid="31004" number="4" />
                <HEAT heatid="31005" number="5" />
                <HEAT heatid="31006" number="6" />
                <HEAT heatid="31007" number="7" />
                <HEAT heatid="31008" number="8" />
                <HEAT heatid="31009" number="9" />
                <HEAT heatid="31010" number="10" />
                <HEAT heatid="31011" number="11" />
                <HEAT heatid="31012" number="12" />
                <HEAT heatid="31013" number="13" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="3" resultid="26" />
                    <RANKING place="4" resultid="335" />
                    <RANKING place="7" resultid="350" />
                    <RANKING place="1" resultid="368" />
                    <RANKING place="6" resultid="1034" />
                    <RANKING place="5" resultid="1247" />
                    <RANKING place="2" resultid="1667" />
                    <RANKING place="8" resultid="1736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="6" resultid="65" />
                    <RANKING place="4" resultid="324" />
                    <RANKING place="1" resultid="604" />
                    <RANKING place="5" resultid="662" />
                    <RANKING place="2" resultid="874" />
                    <RANKING place="3" resultid="1086" />
                    <RANKING place="7" resultid="1122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="9" resultid="74" />
                    <RANKING place="13" resultid="164" />
                    <RANKING place="6" resultid="185" />
                    <RANKING place="2" resultid="194" />
                    <RANKING place="12" resultid="204" />
                    <RANKING place="8" resultid="597" />
                    <RANKING place="11" resultid="837" />
                    <RANKING place="16" resultid="943" />
                    <RANKING place="18" resultid="1107" />
                    <RANKING place="19" resultid="1111" />
                    <RANKING place="15" resultid="1128" />
                    <RANKING place="5" resultid="1190" />
                    <RANKING place="10" resultid="1195" />
                    <RANKING place="3" resultid="1204" />
                    <RANKING place="14" resultid="1210" />
                    <RANKING place="4" resultid="1224" />
                    <RANKING place="1" resultid="1236" />
                    <RANKING place="20" resultid="1686" />
                    <RANKING place="17" resultid="1715" />
                    <RANKING place="7" resultid="1848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="1" resultid="420" />
                    <RANKING place="2" resultid="1115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="170" />
                    <RANKING place="5" resultid="825" />
                    <RANKING place="6" resultid="863" />
                    <RANKING place="3" resultid="902" />
                    <RANKING place="7" resultid="967" />
                    <RANKING place="1" resultid="1699" />
                    <RANKING place="2" resultid="1842" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="32" number="30" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="32000" number="0" />
                <HEAT heatid="32001" number="1" />
                <HEAT heatid="32002" number="2" />
                <HEAT heatid="32003" number="3" />
                <HEAT heatid="32004" number="4" />
                <HEAT heatid="32005" number="5" />
                <HEAT heatid="32006" number="6" />
                <HEAT heatid="32007" number="7" />
                <HEAT heatid="32008" number="8" />
                <HEAT heatid="32009" number="9" />
                <HEAT heatid="32010" number="10" />
                <HEAT heatid="32011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="2" resultid="70" />
                    <RANKING place="1" resultid="229" />
                    <RANKING place="4" resultid="474" />
                    <RANKING place="10" resultid="738" />
                    <RANKING place="7" resultid="890" />
                    <RANKING place="9" resultid="1276" />
                    <RANKING place="3" resultid="1641" />
                    <RANKING place="6" resultid="1778" />
                    <RANKING place="8" resultid="1889" />
                    <RANKING place="5" resultid="1941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="14" resultid="154" />
                    <RANKING place="2" resultid="180" />
                    <RANKING place="12" resultid="199" />
                    <RANKING place="7" resultid="224" />
                    <RANKING place="5" resultid="279" />
                    <RANKING place="17" resultid="345" />
                    <RANKING place="3" resultid="611" />
                    <RANKING place="6" resultid="679" />
                    <RANKING place="11" resultid="761" />
                    <RANKING place="10" resultid="1004" />
                    <RANKING place="13" resultid="1079" />
                    <RANKING place="9" resultid="1176" />
                    <RANKING place="8" resultid="1256" />
                    <RANKING place="1" resultid="1280" />
                    <RANKING place="16" resultid="1496" />
                    <RANKING place="15" resultid="1678" />
                    <RANKING place="18" resultid="1784" />
                    <RANKING place="4" resultid="1836" />
                    <RANKING place="19" resultid="1952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="4" resultid="79" />
                    <RANKING place="7" resultid="395" />
                    <RANKING place="5" resultid="634" />
                    <RANKING place="1" resultid="1092" />
                    <RANKING place="2" resultid="1270" />
                    <RANKING place="3" resultid="1482" />
                    <RANKING place="6" resultid="1822" />
                    <RANKING place="8" resultid="1829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="47" />
                    <RANKING place="2" resultid="657" />
                    <RANKING place="3" resultid="973" />
                    <RANKING place="1" resultid="1171" />
                    <RANKING place="5" resultid="1922" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="33" number="31" gender="F" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="33000" number="0" />
                <HEAT heatid="33001" number="1" />
                <HEAT heatid="33002" number="2" />
                <HEAT heatid="33003" number="3" />
                <HEAT heatid="33004" number="4" />
                <HEAT heatid="33005" number="5" />
                <HEAT heatid="33006" number="6" />
                <HEAT heatid="33007" number="7" />
                <HEAT heatid="33008" number="8" />
                <HEAT heatid="33009" number="9" />
                <HEAT heatid="33010" number="10" />
                <HEAT heatid="33011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="11" resultid="27" />
                    <RANKING place="5" resultid="30" />
                    <RANKING place="7" resultid="42" />
                    <RANKING place="10" resultid="351" />
                    <RANKING place="3" resultid="369" />
                    <RANKING place="8" resultid="571" />
                    <RANKING place="2" resultid="925" />
                    <RANKING place="1" resultid="1010" />
                    <RANKING place="4" resultid="1019" />
                    <RANKING place="9" resultid="1074" />
                    <RANKING place="6" resultid="1248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="10" resultid="66" />
                    <RANKING place="7" resultid="325" />
                    <RANKING place="2" resultid="404" />
                    <RANKING place="8" resultid="466" />
                    <RANKING place="11" resultid="663" />
                    <RANKING place="6" resultid="743" />
                    <RANKING place="1" resultid="875" />
                    <RANKING place="4" resultid="1029" />
                    <RANKING place="3" resultid="1087" />
                    <RANKING place="9" resultid="1558" />
                    <RANKING place="5" resultid="1931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="75" />
                    <RANKING place="6" resultid="165" />
                    <RANKING place="2" resultid="598" />
                    <RANKING place="5" resultid="944" />
                    <RANKING place="7" resultid="1212" />
                    <RANKING place="8" resultid="1716" />
                    <RANKING place="4" resultid="1849" />
                    <RANKING place="9" resultid="1860" />
                    <RANKING place="1" resultid="1874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="1" resultid="144" />
                    <RANKING place="3" resultid="754" />
                    <RANKING place="4" resultid="913" />
                    <RANKING place="2" resultid="1229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="150" />
                    <RANKING place="2" resultid="903" />
                    <RANKING place="4" resultid="968" />
                    <RANKING place="3" resultid="1586" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="34" number="32" gender="M" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="34000" number="0" />
                <HEAT heatid="34001" number="1" />
                <HEAT heatid="34002" number="2" />
                <HEAT heatid="34003" number="3" />
                <HEAT heatid="34004" number="4" />
                <HEAT heatid="34005" number="5" />
                <HEAT heatid="34006" number="6" />
                <HEAT heatid="34007" number="7" />
                <HEAT heatid="34008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="5" resultid="39" />
                    <RANKING place="2" resultid="950" />
                    <RANKING place="1" resultid="1642" />
                    <RANKING place="4" resultid="1779" />
                    <RANKING place="3" resultid="1942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="4" resultid="220" />
                    <RANKING place="9" resultid="400" />
                    <RANKING place="12" resultid="456" />
                    <RANKING place="3" resultid="612" />
                    <RANKING place="10" resultid="1005" />
                    <RANKING place="7" resultid="1065" />
                    <RANKING place="8" resultid="1080" />
                    <RANKING place="1" resultid="1265" />
                    <RANKING place="11" resultid="1497" />
                    <RANKING place="5" resultid="1508" />
                    <RANKING place="6" resultid="1679" />
                    <RANKING place="13" resultid="1785" />
                    <RANKING place="2" resultid="1837" />
                    <RANKING place="14" resultid="1954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="3" resultid="80" />
                    <RANKING place="7" resultid="408" />
                    <RANKING place="4" resultid="635" />
                    <RANKING place="1" resultid="853" />
                    <RANKING place="6" resultid="1479" />
                    <RANKING place="5" resultid="1823" />
                    <RANKING place="2" resultid="1917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="382" />
                    <RANKING place="3" resultid="658" />
                    <RANKING place="5" resultid="897" />
                    <RANKING place="1" resultid="932" />
                    <RANKING place="4" resultid="1260" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="35" number="33" gender="F" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="35001" number="1" />
                <HEAT heatid="35002" number="2" />
                <HEAT heatid="35003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="54" />
                    <RANKING place="5" resultid="186" />
                    <RANKING place="8" resultid="370" />
                    <RANKING place="6" resultid="417" />
                    <RANKING place="9" resultid="914" />
                    <RANKING place="7" resultid="926" />
                    <RANKING place="4" resultid="1191" />
                    <RANKING place="1" resultid="1205" />
                    <RANKING place="3" resultid="1225" />
                    <RANKING place="11" resultid="1737" />
                    <RANKING place="10" resultid="1795" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="36" number="34" gender="M" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="36001" number="1" />
                <HEAT heatid="36002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="383" />
                    <RANKING place="6" resultid="428" />
                    <RANKING place="5" resultid="891" />
                    <RANKING place="3" resultid="1059" />
                    <RANKING place="1" resultid="1172" />
                    <RANKING place="2" resultid="1286" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="37" number="35" gender="F" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="37000" number="0" />
                <HEAT heatid="37001" number="1" />
                <HEAT heatid="37002" number="2" />
                <HEAT heatid="37003" number="3" />
                <HEAT heatid="37004" number="4" />
                <HEAT heatid="37005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="12" resultid="63" />
                    <RANKING place="1" resultid="145" />
                    <RANKING place="3" resultid="171" />
                    <RANKING place="7" resultid="190" />
                    <RANKING place="11" resultid="205" />
                    <RANKING place="9" resultid="257" />
                    <RANKING place="14" resultid="572" />
                    <RANKING place="17" resultid="1075" />
                    <RANKING place="16" resultid="1112" />
                    <RANKING place="3" resultid="1185" />
                    <RANKING place="8" resultid="1196" />
                    <RANKING place="6" resultid="1199" />
                    <RANKING place="2" resultid="1230" />
                    <RANKING place="13" resultid="1696" />
                    <RANKING place="15" resultid="1761" />
                    <RANKING place="18" resultid="1770" />
                    <RANKING place="10" resultid="1870" />
                    <RANKING place="5" resultid="1935" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="38" number="36" gender="M" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="38001" number="1" />
                <HEAT heatid="38002" number="2" />
                <HEAT heatid="38003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="10" resultid="18" />
                    <RANKING place="9" resultid="24" />
                    <RANKING place="4" resultid="71" />
                    <RANKING place="6" resultid="376" />
                    <RANKING place="8" resultid="409" />
                    <RANKING place="7" resultid="475" />
                    <RANKING place="2" resultid="680" />
                    <RANKING place="3" resultid="1177" />
                    <RANKING place="1" resultid="1271" />
                    <RANKING place="5" resultid="1680" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="39" number="37" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="39001" number="1" />
                <HEAT heatid="39002" number="2" />
                <HEAT heatid="39003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Jahrgänge 2013 und älter">
                  <RANKINGS>
                    <RANKING place="6" resultid="313" />
                    <RANKING place="4" resultid="497" />
                    <RANKING place="5" resultid="785" />
                    <RANKING place="3" resultid="994" />
                    <RANKING place="2" resultid="1470" />
                    <RANKING place="1" resultid="1616" />
                    <RANKING place="8" resultid="1622" />
                    <RANKING place="7" resultid="1948" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="40" number="38" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="40001" number="1" />
                <HEAT heatid="40002" number="2" />
                <HEAT heatid="40003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Jahrgänge 2013 und älter">
                  <RANKINGS>
                    <RANKING place="5" resultid="311" />
                    <RANKING place="2" resultid="498" />
                    <RANKING place="3" resultid="783" />
                    <RANKING place="6" resultid="996" />
                    <RANKING place="4" resultid="1474" />
                    <RANKING place="9" resultid="1476" />
                    <RANKING place="1" resultid="1614" />
                    <RANKING place="8" resultid="1620" />
                    <RANKING place="7" resultid="1946" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="4" date="2023-12-10" daytime="13:15">
          <EVENTS>
            <EVENT eventid="41" number="39" gender="F" round="PRE">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="41000" number="0" />
                <HEAT heatid="41001" number="1" />
                <HEAT heatid="41002" number="2" />
                <HEAT heatid="41003" number="3" />
                <HEAT heatid="41004" number="4" />
                <HEAT heatid="41005" number="5" />
                <HEAT heatid="41006" number="6" />
                <HEAT heatid="41007" number="7" />
                <HEAT heatid="41008" number="8" />
                <HEAT heatid="41009" number="9" />
                <HEAT heatid="41010" number="10" />
                <HEAT heatid="41011" number="11" />
                <HEAT heatid="41012" number="12" />
                <HEAT heatid="41013" number="13" />
                <HEAT heatid="41014" number="14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="7" resultid="336" />
                    <RANKING place="5" resultid="352" />
                    <RANKING place="1" resultid="371" />
                    <RANKING place="3" resultid="927" />
                    <RANKING place="2" resultid="1020" />
                    <RANKING place="6" resultid="1249" />
                    <RANKING place="4" resultid="1668" />
                    <RANKING place="8" resultid="1738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="4" resultid="326" />
                    <RANKING place="3" resultid="405" />
                    <RANKING place="9" resultid="467" />
                    <RANKING place="13" resultid="507" />
                    <RANKING place="2" resultid="605" />
                    <RANKING place="10" resultid="664" />
                    <RANKING place="5" resultid="744" />
                    <RANKING place="1" resultid="876" />
                    <RANKING place="7" resultid="1030" />
                    <RANKING place="12" resultid="1039" />
                    <RANKING place="6" resultid="1088" />
                    <RANKING place="14" resultid="1123" />
                    <RANKING place="11" resultid="1559" />
                    <RANKING place="8" resultid="1932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="6" resultid="76" />
                    <RANKING place="11" resultid="166" />
                    <RANKING place="2" resultid="195" />
                    <RANKING place="3" resultid="268" />
                    <RANKING place="7" resultid="599" />
                    <RANKING place="4" resultid="669" />
                    <RANKING place="8" resultid="945" />
                    <RANKING place="9" resultid="1129" />
                    <RANKING place="1" resultid="1243" />
                    <RANKING place="12" resultid="1687" />
                    <RANKING place="10" resultid="1850" />
                    <RANKING place="5" resultid="1875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="1" resultid="55" />
                    <RANKING place="4" resultid="146" />
                    <RANKING place="2" resultid="421" />
                    <RANKING place="5" resultid="755" />
                    <RANKING place="3" resultid="1116" />
                    <RANKING place="6" resultid="1231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="151" />
                    <RANKING place="9" resultid="172" />
                    <RANKING place="8" resultid="826" />
                    <RANKING place="5" resultid="904" />
                    <RANKING place="6" resultid="969" />
                    <RANKING place="7" resultid="1587" />
                    <RANKING place="10" resultid="1700" />
                    <RANKING place="1" resultid="1809" />
                    <RANKING place="3" resultid="1843" />
                    <RANKING place="4" resultid="1936" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="42" number="40" gender="M" round="PRE">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="42000" number="0" />
                <HEAT heatid="42001" number="1" />
                <HEAT heatid="42002" number="2" />
                <HEAT heatid="42003" number="3" />
                <HEAT heatid="42004" number="4" />
                <HEAT heatid="42005" number="5" />
                <HEAT heatid="42006" number="6" />
                <HEAT heatid="42007" number="7" />
                <HEAT heatid="42008" number="8" />
                <HEAT heatid="42009" number="9" />
                <HEAT heatid="42010" number="10" />
                <HEAT heatid="42011" number="11" />
                <HEAT heatid="42012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="3" resultid="377" />
                    <RANKING place="2" resultid="951" />
                    <RANKING place="1" resultid="1643" />
                    <RANKING place="5" resultid="1891" />
                    <RANKING place="4" resultid="1943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="181" />
                    <RANKING place="7" resultid="225" />
                    <RANKING place="4" resultid="280" />
                    <RANKING place="17" resultid="346" />
                    <RANKING place="8" resultid="401" />
                    <RANKING place="10" resultid="457" />
                    <RANKING place="2" resultid="613" />
                    <RANKING place="9" resultid="681" />
                    <RANKING place="11" resultid="762" />
                    <RANKING place="14" resultid="1006" />
                    <RANKING place="13" resultid="1066" />
                    <RANKING place="15" resultid="1081" />
                    <RANKING place="5" resultid="1178" />
                    <RANKING place="6" resultid="1257" />
                    <RANKING place="1" resultid="1281" />
                    <RANKING place="16" resultid="1498" />
                    <RANKING place="12" resultid="1681" />
                    <RANKING place="18" resultid="1953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="4" resultid="81" />
                    <RANKING place="5" resultid="396" />
                    <RANKING place="3" resultid="636" />
                    <RANKING place="1" resultid="854" />
                    <RANKING place="1" resultid="1093" />
                    <RANKING place="9" resultid="1272" />
                    <RANKING place="5" resultid="1287" />
                    <RANKING place="8" resultid="1480" />
                    <RANKING place="10" resultid="1824" />
                    <RANKING place="11" resultid="1830" />
                    <RANKING place="7" resultid="1918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="86" />
                    <RANKING place="5" resultid="366" />
                    <RANKING place="8" resultid="384" />
                    <RANKING place="7" resultid="659" />
                    <RANKING place="6" resultid="898" />
                    <RANKING place="4" resultid="933" />
                    <RANKING place="9" resultid="974" />
                    <RANKING place="11" resultid="1083" />
                    <RANKING place="3" resultid="1173" />
                    <RANKING place="1" resultid="1813" />
                    <RANKING place="10" resultid="1923" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="43" number="41" gender="F" round="PRE">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="43000" number="0" />
                <HEAT heatid="43001" number="1" />
                <HEAT heatid="43002" number="2" />
                <HEAT heatid="43003" number="3" />
                <HEAT heatid="43004" number="4" />
                <HEAT heatid="43005" number="5" />
                <HEAT heatid="43006" number="6" />
                <HEAT heatid="43007" number="7" />
                <HEAT heatid="43008" number="8" />
                <HEAT heatid="43009" number="9" />
                <HEAT heatid="43010" number="10" />
                <HEAT heatid="43011" number="11" />
                <HEAT heatid="43012" number="12" />
                <HEAT heatid="43013" number="13" />
                <HEAT heatid="43014" number="14" />
                <HEAT heatid="43015" number="15" />
                <HEAT heatid="43016" number="16" />
                <HEAT heatid="43017" number="17" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="6" resultid="28" />
                    <RANKING place="5" resultid="337" />
                    <RANKING place="11" resultid="353" />
                    <RANKING place="2" resultid="372" />
                    <RANKING place="8" resultid="573" />
                    <RANKING place="1" resultid="1011" />
                    <RANKING place="3" resultid="1021" />
                    <RANKING place="9" resultid="1036" />
                    <RANKING place="10" resultid="1076" />
                    <RANKING place="7" resultid="1250" />
                    <RANKING place="4" resultid="1669" />
                    <RANKING place="12" resultid="1739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="10" resultid="67" />
                    <RANKING place="4" resultid="327" />
                    <RANKING place="6" resultid="406" />
                    <RANKING place="11" resultid="468" />
                    <RANKING place="12" resultid="508" />
                    <RANKING place="2" resultid="606" />
                    <RANKING place="9" resultid="665" />
                    <RANKING place="1" resultid="877" />
                    <RANKING place="7" resultid="1031" />
                    <RANKING place="3" resultid="1089" />
                    <RANKING place="13" resultid="1124" />
                    <RANKING place="5" resultid="1560" />
                    <RANKING place="8" resultid="1933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="15" resultid="77" />
                    <RANKING place="17" resultid="167" />
                    <RANKING place="8" resultid="187" />
                    <RANKING place="2" resultid="196" />
                    <RANKING place="16" resultid="206" />
                    <RANKING place="4" resultid="269" />
                    <RANKING place="5" resultid="670" />
                    <RANKING place="11" resultid="781" />
                    <RANKING place="10" resultid="838" />
                    <RANKING place="18" resultid="946" />
                    <RANKING place="22" resultid="1108" />
                    <RANKING place="21" resultid="1130" />
                    <RANKING place="6" resultid="1181" />
                    <RANKING place="14" resultid="1186" />
                    <RANKING place="9" resultid="1192" />
                    <RANKING place="3" resultid="1206" />
                    <RANKING place="20" resultid="1211" />
                    <RANKING place="7" resultid="1226" />
                    <RANKING place="1" resultid="1237" />
                    <RANKING place="24" resultid="1688" />
                    <RANKING place="19" resultid="1717" />
                    <RANKING place="13" resultid="1851" />
                    <RANKING place="23" resultid="1861" />
                    <RANKING place="12" resultid="1876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="1" resultid="56" />
                    <RANKING place="2" resultid="422" />
                    <RANKING place="5" resultid="915" />
                    <RANKING place="4" resultid="1117" />
                    <RANKING place="3" resultid="1232" />
                    <RANKING place="6" resultid="1908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="152" />
                    <RANKING place="8" resultid="827" />
                    <RANKING place="9" resultid="864" />
                    <RANKING place="4" resultid="905" />
                    <RANKING place="6" resultid="1588" />
                    <RANKING place="7" resultid="1701" />
                    <RANKING place="1" resultid="1810" />
                    <RANKING place="3" resultid="1844" />
                    <RANKING place="5" resultid="1937" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="44" number="42" gender="M" round="PRE">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="44000" number="0" />
                <HEAT heatid="44001" number="1" />
                <HEAT heatid="44002" number="2" />
                <HEAT heatid="44003" number="3" />
                <HEAT heatid="44004" number="4" />
                <HEAT heatid="44005" number="5" />
                <HEAT heatid="44006" number="6" />
                <HEAT heatid="44007" number="7" />
                <HEAT heatid="44008" number="8" />
                <HEAT heatid="44009" number="9" />
                <HEAT heatid="44010" number="10" />
                <HEAT heatid="44011" number="11" />
                <HEAT heatid="44012" number="12" />
                <HEAT heatid="44013" number="13" />
                <HEAT heatid="44014" number="14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="2" resultid="72" />
                    <RANKING place="6" resultid="378" />
                    <RANKING place="3" resultid="476" />
                    <RANKING place="10" resultid="739" />
                    <RANKING place="8" resultid="892" />
                    <RANKING place="7" resultid="1277" />
                    <RANKING place="1" resultid="1644" />
                    <RANKING place="4" resultid="1781" />
                    <RANKING place="9" resultid="1892" />
                    <RANKING place="5" resultid="1944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="17" resultid="155" />
                    <RANKING place="2" resultid="182" />
                    <RANKING place="18" resultid="200" />
                    <RANKING place="8" resultid="221" />
                    <RANKING place="9" resultid="226" />
                    <RANKING place="20" resultid="347" />
                    <RANKING place="10" resultid="402" />
                    <RANKING place="15" resultid="458" />
                    <RANKING place="4" resultid="614" />
                    <RANKING place="7" resultid="682" />
                    <RANKING place="12" resultid="763" />
                    <RANKING place="13" resultid="1007" />
                    <RANKING place="11" resultid="1082" />
                    <RANKING place="1" resultid="1266" />
                    <RANKING place="3" resultid="1282" />
                    <RANKING place="19" resultid="1499" />
                    <RANKING place="6" resultid="1509" />
                    <RANKING place="15" resultid="1682" />
                    <RANKING place="14" resultid="1786" />
                    <RANKING place="5" resultid="1838" />
                    <RANKING place="21" resultid="1955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="5" resultid="82" />
                    <RANKING place="7" resultid="397" />
                    <RANKING place="11" resultid="410" />
                    <RANKING place="1" resultid="637" />
                    <RANKING place="2" resultid="855" />
                    <RANKING place="10" resultid="1060" />
                    <RANKING place="4" resultid="1094" />
                    <RANKING place="6" resultid="1288" />
                    <RANKING place="3" resultid="1483" />
                    <RANKING place="8" resultid="1825" />
                    <RANKING place="12" resultid="1831" />
                    <RANKING place="9" resultid="1919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="87" />
                    <RANKING place="7" resultid="660" />
                    <RANKING place="4" resultid="934" />
                    <RANKING place="6" resultid="975" />
                    <RANKING place="9" resultid="1084" />
                    <RANKING place="3" resultid="1174" />
                    <RANKING place="5" resultid="1261" />
                    <RANKING place="1" resultid="1814" />
                    <RANKING place="8" resultid="1924" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="45" number="43" gender="F" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="45000" number="0" />
                <HEAT heatid="45001" number="1" />
                <HEAT heatid="45002" number="2" />
                <HEAT heatid="45003" number="3" />
                <HEAT heatid="45004" number="4" />
                <HEAT heatid="45005" number="5" />
                <HEAT heatid="45006" number="6" />
                <HEAT heatid="45007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="1" resultid="31" />
                    <RANKING place="2" resultid="574" />
                    <RANKING place="4" resultid="1037" />
                    <RANKING place="3" resultid="1077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="2" resultid="745" />
                    <RANKING place="3" resultid="1041" />
                    <RANKING place="1" resultid="1934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="6" resultid="207" />
                    <RANKING place="5" resultid="258" />
                    <RANKING place="7" resultid="1113" />
                    <RANKING place="1" resultid="1182" />
                    <RANKING place="4" resultid="1187" />
                    <RANKING place="2" resultid="1197" />
                    <RANKING place="3" resultid="1200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="2" resultid="147" />
                    <RANKING place="3" resultid="191" />
                    <RANKING place="1" resultid="1233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="173" />
                    <RANKING place="2" resultid="828" />
                    <RANKING place="3" resultid="865" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="46" number="44" gender="M" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="46000" number="0" />
                <HEAT heatid="46001" number="1" />
                <HEAT heatid="46002" number="2" />
                <HEAT heatid="46003" number="3" />
                <HEAT heatid="46004" number="4" />
                <HEAT heatid="46005" number="5" />
                <HEAT heatid="46006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="1" resultid="73" />
                    <RANKING place="4" resultid="379" />
                    <RANKING place="2" resultid="477" />
                    <RANKING place="5" resultid="740" />
                    <RANKING place="3" resultid="1645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="3" resultid="201" />
                    <RANKING place="1" resultid="683" />
                    <RANKING place="2" resultid="1067" />
                    <RANKING place="5" resultid="1500" />
                    <RANKING place="7" resultid="1510" />
                    <RANKING place="4" resultid="1683" />
                    <RANKING place="6" resultid="1787" />
                    <RANKING place="8" resultid="1956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="4" resultid="411" />
                    <RANKING place="3" resultid="1061" />
                    <RANKING place="1" resultid="1273" />
                    <RANKING place="5" resultid="1832" />
                    <RANKING place="2" resultid="1920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="385" />
                    <RANKING place="2" resultid="899" />
                    <RANKING place="3" resultid="976" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="47" number="45" gender="F" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="47001" number="1" />
                <HEAT heatid="47002" number="2" />
                <HEAT heatid="47003" number="3" />
                <HEAT heatid="47004" number="4" />
                <HEAT heatid="47005" number="5" />
                <HEAT heatid="47006" number="6" />
                <HEAT heatid="47007" number="7" />
                <HEAT heatid="47008" number="8" />
                <HEAT heatid="47009" number="9" />
                <HEAT heatid="47010" number="10" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="6" resultid="43" />
                    <RANKING place="3" resultid="373" />
                    <RANKING place="2" resultid="928" />
                    <RANKING place="1" resultid="1012" />
                    <RANKING place="4" resultid="1022" />
                    <RANKING place="5" resultid="1670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="2" resultid="607" />
                    <RANKING place="6" resultid="666" />
                    <RANKING place="3" resultid="746" />
                    <RANKING place="1" resultid="878" />
                    <RANKING place="4" resultid="1032" />
                    <RANKING place="5" resultid="1561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="11" resultid="168" />
                    <RANKING place="6" resultid="600" />
                    <RANKING place="5" resultid="782" />
                    <RANKING place="10" resultid="839" />
                    <RANKING place="9" resultid="947" />
                    <RANKING place="12" resultid="1109" />
                    <RANKING place="7" resultid="1188" />
                    <RANKING place="4" resultid="1193" />
                    <RANKING place="1" resultid="1207" />
                    <RANKING place="14" resultid="1208" />
                    <RANKING place="3" resultid="1227" />
                    <RANKING place="2" resultid="1238" />
                    <RANKING place="16" resultid="1689" />
                    <RANKING place="13" resultid="1718" />
                    <RANKING place="8" resultid="1852" />
                    <RANKING place="15" resultid="1862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="1" resultid="57" />
                    <RANKING place="2" resultid="1118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="970" />
                    <RANKING place="3" resultid="1589" />
                    <RANKING place="1" resultid="1702" />
                    <RANKING place="2" resultid="1845" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="48" number="46" gender="M" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="48001" number="1" />
                <HEAT heatid="48002" number="2" />
                <HEAT heatid="48003" number="3" />
                <HEAT heatid="48004" number="4" />
                <HEAT heatid="48005" number="5" />
                <HEAT heatid="48006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="3" resultid="893" />
                    <RANKING place="2" resultid="952" />
                    <RANKING place="4" resultid="1782" />
                    <RANKING place="5" resultid="1893" />
                    <RANKING place="1" resultid="1945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="7" resultid="156" />
                    <RANKING place="3" resultid="281" />
                    <RANKING place="6" resultid="348" />
                    <RANKING place="5" resultid="615" />
                    <RANKING place="2" resultid="1267" />
                    <RANKING place="4" resultid="1839" />
                    <RANKING place="1" resultid="1939" />
                    <RANKING place="8" resultid="1957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="2" resultid="638" />
                    <RANKING place="3" resultid="1062" />
                    <RANKING place="1" resultid="1289" />
                    <RANKING place="4" resultid="1484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="48" />
                    <RANKING place="3" resultid="661" />
                    <RANKING place="5" resultid="977" />
                    <RANKING place="1" resultid="1175" />
                    <RANKING place="2" resultid="1262" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="49" number="47" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="200" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="49001" number="1" />
                <HEAT heatid="49002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="192" />
                    <RANKING place="5" resultid="756" />
                    <RANKING place="4" resultid="1201" />
                    <RANKING place="2" resultid="1244" />
                    <RANKING place="6" resultid="1251" />
                    <RANKING place="1" resultid="1938" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="50" number="48" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="50001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="11" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="230" />
                    <RANKING place="1" resultid="1283" />
                    <RANKING place="3" resultid="1646" />
                    <RANKING place="4" resultid="1833" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="51" number="49" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="51001" number="1" />
                <HEAT heatid="51002" number="2" />
                <HEAT heatid="51003" number="3" />
                <HEAT heatid="51004" number="4" />
                <HEAT heatid="51005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="9" resultid="64" />
                    <RANKING place="5" resultid="68" />
                    <RANKING place="3" resultid="188" />
                    <RANKING place="2" resultid="197" />
                    <RANKING place="8" resultid="328" />
                    <RANKING place="12" resultid="338" />
                    <RANKING place="7" resultid="418" />
                    <RANKING place="13" resultid="1125" />
                    <RANKING place="1" resultid="1239" />
                    <RANKING place="14" resultid="1697" />
                    <RANKING place="16" resultid="1740" />
                    <RANKING place="10" resultid="1762" />
                    <RANKING place="15" resultid="1771" />
                    <RANKING place="4" resultid="1846" />
                    <RANKING place="11" resultid="1871" />
                    <RANKING place="6" resultid="1877" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="52" number="50" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="52001" number="1" />
                <HEAT heatid="52002" number="2" />
                <HEAT heatid="52003" number="3" />
                <HEAT heatid="52004" number="4" />
                <HEAT heatid="52005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="12" resultid="19" />
                    <RANKING place="13" resultid="25" />
                    <RANKING place="3" resultid="83" />
                    <RANKING place="10" resultid="157" />
                    <RANKING place="4" resultid="183" />
                    <RANKING place="5" resultid="222" />
                    <RANKING place="8" resultid="227" />
                    <RANKING place="6" resultid="231" />
                    <RANKING place="11" resultid="429" />
                    <RANKING place="9" resultid="764" />
                    <RANKING place="1" resultid="856" />
                    <RANKING place="15" resultid="1278" />
                    <RANKING place="2" resultid="1284" />
                    <RANKING place="7" resultid="1826" />
                    <RANKING place="14" resultid="1894" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="53" number="51" gender="F" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="53001" number="1" />
                <HEAT heatid="53002" number="2" />
                <HEAT heatid="53003" number="3" />
                <HEAT heatid="53004" number="4" />
                <HEAT heatid="53005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="13" agemin="13" name="Jahrgang 2010">
                  <RANKINGS>
                    <RANKING place="2" resultid="354" />
                    <RANKING place="1" resultid="1671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009" />
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="2" resultid="78" />
                    <RANKING place="4" resultid="259" />
                    <RANKING place="3" resultid="601" />
                    <RANKING place="1" resultid="1245" />
                    <RANKING place="5" resultid="1863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="2" resultid="58" />
                    <RANKING place="1" resultid="423" />
                    <RANKING place="3" resultid="757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="906" />
                    <RANKING place="2" resultid="971" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="54" number="52" gender="M" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="54001" number="1" />
                <HEAT heatid="54002" number="2" />
                <HEAT heatid="54003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="14" name="Jahrgang 2009">
                  <RANKINGS>
                    <RANKING place="3" resultid="40" />
                    <RANKING place="2" resultid="953" />
                    <RANKING place="1" resultid="1647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="16" agemin="15" name="Jahrgänge 2007/2008">
                  <RANKINGS>
                    <RANKING place="2" resultid="202" />
                    <RANKING place="1" resultid="684" />
                    <RANKING place="4" resultid="1684" />
                    <RANKING place="3" resultid="1788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="17" name="Jahrgänge 2005/2006">
                  <RANKINGS>
                    <RANKING place="1" resultid="857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="Jahrgänge 2004 und älter">
                  <RANKINGS>
                    <RANKING place="2" resultid="386" />
                    <RANKING place="1" resultid="1120" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="55" number="123" gender="F" round="FIN">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="55001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2037" />
                    <RANKING place="2" resultid="2038" />
                    <RANKING place="4" resultid="2039" />
                    <RANKING place="3" resultid="2040" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="56" number="223" gender="F" round="FIN">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="56001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="13" name="2010 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2041" />
                    <RANKING place="4" resultid="2042" />
                    <RANKING place="2" resultid="2043" />
                    <RANKING place="3" resultid="2044" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="16" agemin="13" name="Juniorenwertung" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="57" number="124" gender="M" round="FIN">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="57001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2045" />
                    <RANKING place="4" resultid="2046" />
                    <RANKING place="3" resultid="2047" />
                    <RANKING place="2" resultid="2048" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="58" number="224" gender="M" round="FIN">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="58001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="14" name="2009 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2049" />
                    <RANKING place="2" resultid="2050" />
                    <RANKING place="3" resultid="2051" />
                    <RANKING place="4" resultid="2052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Juniorenwertung" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="59" number="125" gender="F" round="FIN">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="59001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="2053" />
                    <RANKING place="3" resultid="2054" />
                    <RANKING place="4" resultid="2055" />
                    <RANKING place="5" resultid="2056" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="60" number="225" gender="F" round="FIN">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="60001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="13" name="2010 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2057" />
                    <RANKING place="4" resultid="2058" />
                    <RANKING place="3" resultid="2059" />
                    <RANKING place="2" resultid="2060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2058" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="61" number="126" gender="M" round="FIN">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="61000" number="0" />
                <HEAT heatid="61001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="2062" />
                    <RANKING place="2" resultid="2063" />
                    <RANKING place="4" resultid="2064" />
                    <RANKING place="5" resultid="2065" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="62" number="226" gender="M" round="FIN">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="62000" number="0" />
                <HEAT heatid="62001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="14" name="2009 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2067" />
                    <RANKING place="2" resultid="2068" />
                    <RANKING place="3" resultid="2069" />
                    <RANKING place="4" resultid="2070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2070" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="63" number="139" gender="F" round="FIN">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="63001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2071" />
                    <RANKING place="2" resultid="2072" />
                    <RANKING place="3" resultid="2073" />
                    <RANKING place="4" resultid="2074" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="64" number="239" gender="F" round="FIN">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="64001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="13" name="2010 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2075" />
                    <RANKING place="2" resultid="2076" />
                    <RANKING place="3" resultid="2077" />
                    <RANKING place="4" resultid="2078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="16" agemin="13" name="Juniorenwertung" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="65" number="140" gender="M" round="FIN">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="65001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="2079" />
                    <RANKING place="4" resultid="2080" />
                    <RANKING place="5" resultid="2081" />
                    <RANKING place="2" resultid="2082" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="66" number="240" gender="M" round="FIN">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="66001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="14" name="2009 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2083" />
                    <RANKING place="2" resultid="2084" />
                    <RANKING place="3" resultid="2085" />
                    <RANKING place="4" resultid="2086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2086" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="67" number="141" gender="F" round="FIN">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="67001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="16" agemin="13" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2087" />
                    <RANKING place="2" resultid="2088" />
                    <RANKING place="4" resultid="2089" />
                    <RANKING place="3" resultid="2090" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="68" number="241" gender="F" round="FIN">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="68001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="13" name="2010 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2091" />
                    <RANKING place="4" resultid="2092" />
                    <RANKING place="2" resultid="2093" />
                    <RANKING place="3" resultid="2094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="16" agemin="13" name="Juniorenwertung" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="69" number="142" gender="M" round="FIN">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="69000" number="0" />
                <HEAT heatid="69001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="17" agemin="12" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="2096" />
                    <RANKING place="3" resultid="2097" />
                    <RANKING place="4" resultid="2098" />
                    <RANKING place="5" resultid="2099" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="70" number="242" gender="M" round="FIN">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="70001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="14" name="2009 und älter">
                  <RANKINGS>
                    <RANKING place="1" resultid="2100" />
                    <RANKING place="2" resultid="2101" />
                    <RANKING place="4" resultid="2102" />
                    <RANKING place="3" resultid="2103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Juniorenwertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2102" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="71" number="53" gender="F" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="71001" number="1" />
                <HEAT heatid="71002" number="2" />
                <HEAT heatid="71003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Jahrgänge 2013 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="499" />
                    <RANKING place="3" resultid="786" />
                    <RANKING place="6" resultid="995" />
                    <RANKING place="1" resultid="1471" />
                    <RANKING place="2" resultid="1617" />
                    <RANKING place="7" resultid="1623" />
                    <RANKING place="8" resultid="1627" />
                    <RANKING place="5" resultid="1949" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="72" number="54" gender="M" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="72001" number="1" />
                <HEAT heatid="72002" number="2" />
                <HEAT heatid="72003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="10" name="Jahrgänge 2013 und älter">
                  <RANKINGS>
                    <RANKING place="4" resultid="500" />
                    <RANKING place="2" resultid="784" />
                    <RANKING place="5" resultid="997" />
                    <RANKING place="1" resultid="1475" />
                    <RANKING place="7" resultid="1477" />
                    <RANKING place="3" resultid="1615" />
                    <RANKING place="8" resultid="1621" />
                    <RANKING place="9" resultid="1626" />
                    <RANKING place="6" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="ATSV Freiberg e.V." nation="GER" region="12" code="3324">
          <ATHLETES>
            <ATHLETE athleteid="325" birthdate="2013-01-01" gender="F" lastname="Brocke" firstname="Fiene" license="445947">
              <RESULTS>
                <RESULT resultid="1489" eventid="1" swimtime="00:01:57.64" lane="3" heatid="1001">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:54.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1490" eventid="3" swimtime="00:00:51.66" lane="3" heatid="3008" />
                <RESULT resultid="1491" eventid="9" swimtime="00:01:51.12" lane="2" heatid="9004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1492" eventid="13" swimtime="00:00:55.33" lane="2" heatid="13002" />
                <RESULT resultid="1493" eventid="17" swimtime="00:00:56.20" lane="2" heatid="17005" />
                <RESULT resultid="1494" eventid="19" swimtime="00:01:44.52" lane="1" heatid="19004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="326" birthdate="2007-01-01" gender="M" lastname="Frisch" firstname="Jonathan" license="384470">
              <RESULTS>
                <RESULT resultid="1495" eventid="28" swimtime="00:00:36.82" lane="4" heatid="28003" />
                <RESULT resultid="1496" eventid="32" swimtime="00:01:08.29" lane="1" heatid="32003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1497" eventid="34" swimtime="00:01:17.55" lane="3" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1498" eventid="42" swimtime="00:00:34.29" lane="1" heatid="42002" />
                <RESULT resultid="1499" eventid="44" swimtime="00:00:30.41" lane="3" heatid="44003" />
                <RESULT resultid="1500" eventid="46" swimtime="00:01:24.83" lane="2" heatid="46002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="327" birthdate="2014-01-01" gender="F" lastname="Grämer" firstname="Stella" license="445949">
              <RESULTS>
                <RESULT resultid="1501" eventid="3" status="DSQ" swimtime="00:00:47.96" lane="4" heatid="3005" comment="Die Sportlerin hat bei der Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt." />
                <RESULT resultid="1502" eventid="7" swimtime="00:00:40.32" lane="3" heatid="7010" />
                <RESULT resultid="1503" eventid="9" swimtime="00:01:46.23" lane="2" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1504" eventid="13" swimtime="00:00:48.84" lane="1" heatid="13007" />
                <RESULT resultid="1505" eventid="15" status="DSQ" swimtime="00:01:45.47" lane="4" heatid="15005" comment="Die Sportlerin hat bei der dritten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1506" eventid="19" swimtime="00:01:35.70" lane="1" heatid="19005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="328" birthdate="2008-01-01" gender="M" lastname="Heinrich" firstname="Tim" license="364363">
              <RESULTS>
                <RESULT resultid="1507" eventid="28" swimtime="00:00:34.29" lane="4" heatid="28007" />
                <RESULT resultid="1508" eventid="34" swimtime="00:01:11.75" lane="4" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1509" eventid="44" swimtime="00:00:26.28" lane="4" heatid="44009" />
                <RESULT resultid="1510" eventid="46" swimtime="00:01:25.54" lane="2" heatid="46001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2061" eventid="61" status="WDR" swimtime="00:00:00.00" lane="0" heatid="61000" />
                <RESULT resultid="2095" eventid="69" status="WDR" swimtime="00:00:00.00" lane="0" heatid="69000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="329" birthdate="2015-01-01" gender="F" lastname="Heinz" firstname="Elizabeth" license="471931">
              <RESULTS>
                <RESULT resultid="1511" eventid="3" status="DSQ" swimtime="00:00:55.81" lane="1" heatid="3006" comment="Die Sportlerin hat bei der Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt." />
                <RESULT resultid="1512" eventid="5" swimtime="00:02:17.46" lane="4" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1513" eventid="7" status="DSQ" swimtime="00:00:49.53" lane="3" heatid="7005" comment="Dier Sportlerin startete vor dem Startsignal" />
                <RESULT resultid="1514" eventid="15" swimtime="00:01:57.13" lane="4" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1515" eventid="17" swimtime="00:00:58.82" lane="4" heatid="17010" />
                <RESULT resultid="1516" eventid="19" swimtime="00:01:54.30" lane="2" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="330" birthdate="2014-01-01" gender="F" lastname="Irmscher" firstname="Nora" license="445948">
              <RESULTS>
                <RESULT resultid="1517" eventid="3" swimtime="00:00:54.67" lane="3" heatid="3005" />
                <RESULT resultid="1518" eventid="7" swimtime="00:00:45.72" lane="1" heatid="7007" />
                <RESULT resultid="1519" eventid="9" swimtime="00:02:00.18" lane="1" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="331" birthdate="2012-01-01" gender="F" lastname="Kaiser" firstname="Zoe" license="431997">
              <RESULTS>
                <RESULT resultid="1520" eventid="1" swimtime="00:01:32.38" lane="1" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1521" eventid="3" swimtime="00:00:42.39" lane="2" heatid="3016" />
                <RESULT resultid="1522" eventid="7" swimtime="00:00:34.18" lane="3" heatid="7015" />
                <RESULT resultid="1523" eventid="13" swimtime="00:00:40.75" lane="2" heatid="13004" />
                <RESULT resultid="1524" eventid="15" swimtime="00:01:32.47" lane="2" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1525" eventid="19" swimtime="00:01:24.39" lane="4" heatid="19010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="332" birthdate="2012-01-01" gender="F" lastname="Michel" firstname="Virsavia" license="434284">
              <RESULTS>
                <RESULT resultid="1526" eventid="3" swimtime="00:00:41.71" lane="4" heatid="3016" />
                <RESULT resultid="1527" eventid="5" swimtime="00:01:42.14" lane="4" heatid="5007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1528" eventid="9" swimtime="00:01:29.82" lane="2" heatid="9009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1529" eventid="13" swimtime="00:00:42.54" lane="3" heatid="13004" />
                <RESULT resultid="1530" eventid="17" swimtime="00:00:45.60" lane="1" heatid="17013" />
                <RESULT resultid="1531" eventid="19" swimtime="00:01:19.82" lane="3" heatid="19010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="333" birthdate="2013-01-01" gender="F" lastname="Müller" firstname="Lara" license="431998">
              <RESULTS>
                <RESULT resultid="1532" eventid="3" swimtime="00:00:58.00" lane="1" heatid="3004" />
                <RESULT resultid="1533" eventid="7" swimtime="00:00:49.27" lane="1" heatid="7006" />
                <RESULT resultid="1534" eventid="9" swimtime="00:02:09.07" lane="2" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1535" eventid="13" swimtime="00:01:00.39" lane="3" heatid="13001" />
                <RESULT resultid="1536" eventid="15" swimtime="00:02:10.17" lane="3" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1537" eventid="19" swimtime="00:01:58.66" lane="3" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="334" birthdate="2013-01-01" gender="M" lastname="Oehme" firstname="Arvid" license="445060">
              <RESULTS>
                <RESULT resultid="1538" eventid="2" swimtime="00:01:45.49" lane="4" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:45.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1539" eventid="8" swimtime="00:00:37.74" lane="4" heatid="8009" />
                <RESULT resultid="1540" eventid="10" swimtime="00:01:34.68" lane="1" heatid="10004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1541" eventid="14" swimtime="00:00:41.26" lane="1" heatid="14006" />
                <RESULT resultid="1542" eventid="18" swimtime="00:00:51.39" lane="2" heatid="18005" />
                <RESULT resultid="1543" eventid="20" swimtime="00:01:28.61" lane="2" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="335" birthdate="2013-01-01" gender="F" lastname="Queck" firstname="Fabienne" license="451852">
              <RESULTS>
                <RESULT resultid="1544" eventid="5" swimtime="00:01:53.22" lane="2" heatid="5003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1545" eventid="7" swimtime="00:00:43.01" lane="2" heatid="7007" />
                <RESULT resultid="1546" eventid="9" swimtime="00:01:51.73" lane="3" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1547" eventid="13" swimtime="00:00:56.30" lane="1" heatid="13002" />
                <RESULT resultid="1548" eventid="17" swimtime="00:00:50.39" lane="4" heatid="17007" />
                <RESULT resultid="1549" eventid="19" swimtime="00:01:41.27" lane="3" heatid="19003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="336" birthdate="2011-01-01" gender="M" lastname="Rülke" firstname="Luca" license="431995">
              <RESULTS>
                <RESULT resultid="1550" eventid="4" swimtime="00:00:50.06" lane="2" heatid="4003" />
                <RESULT resultid="1551" eventid="6" swimtime="00:01:58.16" lane="4" heatid="6004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1552" eventid="8" swimtime="00:00:40.57" lane="3" heatid="8008" />
                <RESULT resultid="1553" eventid="16" swimtime="00:01:47.37" lane="4" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1554" eventid="18" swimtime="00:00:54.00" lane="1" heatid="18004" />
                <RESULT resultid="1555" eventid="20" swimtime="00:01:36.98" lane="3" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="337" birthdate="2009-01-01" gender="F" lastname="Schierz" firstname="Johanna" license="383730">
              <RESULTS>
                <RESULT resultid="1556" eventid="25" status="DSQ" swimtime="00:00:34.48" lane="4" heatid="25010" comment="Vor der Wende führte die Sportlerin in Bauchlage zwei Armzüge aus." />
                <RESULT resultid="1557" eventid="27" swimtime="00:00:43.18" lane="2" heatid="27003" />
                <RESULT resultid="1558" eventid="33" swimtime="00:01:23.01" lane="1" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1559" eventid="41" swimtime="00:00:37.45" lane="2" heatid="41002" />
                <RESULT resultid="1560" eventid="43" swimtime="00:00:30.63" lane="2" heatid="43011" />
                <RESULT resultid="1561" eventid="47" swimtime="00:01:23.95" lane="4" heatid="47005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="338" birthdate="2012-01-01" gender="M" lastname="Schubert" firstname="Fritz" license="422021">
              <RESULTS>
                <RESULT resultid="1562" eventid="4" status="DSQ" swimtime="00:00:41.67" lane="2" heatid="4008" comment="Der Sportler hat bei der Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt." />
                <RESULT resultid="1563" eventid="8" swimtime="00:00:33.44" lane="4" heatid="8018" />
                <RESULT resultid="1564" eventid="10" swimtime="00:01:30.41" lane="2" heatid="10004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1565" eventid="14" swimtime="00:00:41.99" lane="2" heatid="14004" />
                <RESULT resultid="1566" eventid="16" swimtime="00:01:30.48" lane="1" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1567" eventid="20" swimtime="00:01:13.78" lane="3" heatid="20010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="339" birthdate="2012-01-01" gender="M" lastname="Tanneberger" firstname="Arian" license="434981">
              <RESULTS>
                <RESULT resultid="1568" eventid="2" swimtime="00:01:41.88" lane="4" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1569" eventid="6" swimtime="00:01:44.71" lane="4" heatid="6008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1570" eventid="8" swimtime="00:00:33.71" lane="1" heatid="8018" />
                <RESULT resultid="1571" eventid="14" swimtime="00:00:41.13" lane="4" heatid="14009" />
                <RESULT resultid="1572" eventid="18" swimtime="00:00:48.97" lane="2" heatid="18006" />
                <RESULT resultid="1573" eventid="20" swimtime="00:01:18.05" lane="4" heatid="20014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="340" birthdate="2010-01-01" gender="M" lastname="Tanneberger" firstname="Janis" license="407515">
              <RESULTS>
                <RESULT resultid="1574" eventid="4" swimtime="00:00:37.30" lane="3" heatid="4015" />
                <RESULT resultid="1575" eventid="6" swimtime="00:01:37.68" lane="1" heatid="6010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1576" eventid="8" swimtime="00:00:32.87" lane="3" heatid="8014" />
                <RESULT resultid="1577" eventid="14" swimtime="00:00:36.97" lane="4" heatid="14011" />
                <RESULT resultid="1578" eventid="16" swimtime="00:01:24.41" lane="1" heatid="16009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1579" eventid="18" swimtime="00:00:42.70" lane="3" heatid="18013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="341" birthdate="1989-01-01" gender="F" lastname="Weßolowski" firstname="Carolin" license="172726">
              <RESULTS>
                <RESULT resultid="1580" eventid="29" status="WDR" swimtime="00:00:00.00" lane="0" heatid="29000" />
                <RESULT resultid="1581" eventid="33" status="WDR" swimtime="00:00:00.00" lane="0" heatid="33000" />
                <RESULT resultid="1582" eventid="41" status="WDR" swimtime="00:00:00.00" lane="0" heatid="41000" />
                <RESULT resultid="1583" eventid="45" status="WDR" swimtime="00:00:00.00" lane="0" heatid="45000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="342" birthdate="2003-01-01" gender="F" lastname="Wolf" firstname="Leonie" license="242026">
              <RESULTS>
                <RESULT resultid="1584" eventid="25" swimtime="00:00:35.41" lane="4" heatid="25008" />
                <RESULT resultid="1585" eventid="27" swimtime="00:00:40.96" lane="1" heatid="27009" />
                <RESULT resultid="1586" eventid="33" swimtime="00:01:18.08" lane="1" heatid="33011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1587" eventid="41" swimtime="00:00:33.28" lane="3" heatid="41008" />
                <RESULT resultid="1588" eventid="43" swimtime="00:00:30.29" lane="4" heatid="43010" />
                <RESULT resultid="1589" eventid="47" swimtime="00:01:16.92" lane="1" heatid="47010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1488" eventid="11" swimtime="00:02:12.54" lane="2" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:06.11" />
                    <SPLIT distance="150" swimtime="00:01:39.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="340" number="1" />
                    <RELAYPOSITION athleteid="332" number="2" />
                    <RELAYPOSITION athleteid="339" number="3" />
                    <RELAYPOSITION athleteid="338" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Berliner TSC" nation="GER" region="3" code="5650">
          <ATHLETES>
            <ATHLETE athleteid="413" birthdate="2000-01-01" gender="F" lastname="Gränitz" firstname="Hanka" license="292499">
              <RESULTS>
                <RESULT resultid="1935" eventid="37" swimtime="00:02:58.39" lane="4" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                    <SPLIT distance="100" swimtime="00:01:25.79" />
                    <SPLIT distance="150" swimtime="00:02:11.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1936" eventid="41" swimtime="00:00:32.19" lane="3" heatid="41009" />
                <RESULT resultid="1937" eventid="43" swimtime="00:00:29.95" lane="3" heatid="43012" />
                <RESULT resultid="1938" eventid="49" swimtime="00:02:32.83" lane="2" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:50.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="BKS Swim Team Bielawa" nation="POL" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="242" birthdate="2011-01-01" gender="F" lastname="Boczar" firstname="Roksana" license="0">
              <RESULTS>
                <RESULT resultid="1131" eventid="5" swimtime="00:01:32.31" lane="3" heatid="5001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1132" eventid="7" swimtime="00:00:34.39" lane="3" heatid="7013" />
                <RESULT resultid="1133" eventid="17" swimtime="00:00:41.34" lane="1" heatid="17007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="243" birthdate="2011-01-01" gender="F" lastname="Cergier" firstname="Samanta" license="0">
              <RESULTS>
                <RESULT resultid="1134" eventid="5" swimtime="00:01:49.74" lane="2" heatid="5001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1135" eventid="7" swimtime="00:00:40.48" lane="4" heatid="7012" />
                <RESULT resultid="1136" eventid="17" swimtime="00:00:51.26" lane="2" heatid="17006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="244" birthdate="2010-01-01" gender="M" lastname="Ciosek" firstname="Jakub" license="0">
              <RESULTS>
                <RESULT resultid="1137" eventid="8" swimtime="00:00:29.50" lane="1" heatid="8020" />
                <RESULT resultid="1138" eventid="10" swimtime="00:01:19.16" lane="1" heatid="10011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1139" eventid="20" swimtime="00:01:09.93" lane="1" heatid="20016">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="245" birthdate="2013-01-01" gender="M" lastname="Dabrowski" firstname="Leon" license="0">
              <RESULTS>
                <RESULT resultid="1140" eventid="8" swimtime="00:00:49.36" lane="3" heatid="8002" />
                <RESULT resultid="1141" eventid="18" status="DSQ" swimtime="00:00:58.05" lane="4" heatid="18004" comment="Nach dem Start hat der Sportler zwei Tauchzüge ausgeführt." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="246" birthdate="2013-01-01" gender="M" lastname="Denysiewicz" firstname="Piotr" license="0">
              <RESULTS>
                <RESULT resultid="1142" eventid="6" swimtime="00:01:48.30" lane="2" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1143" eventid="8" swimtime="00:00:40.59" lane="3" heatid="8010" />
                <RESULT resultid="1144" eventid="18" swimtime="00:00:50.63" lane="4" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="247" birthdate="2011-01-01" gender="F" lastname="Dziedzic" firstname="Maja" license="0">
              <RESULTS>
                <RESULT resultid="1145" eventid="3" swimtime="00:00:45.44" lane="1" heatid="3001" />
                <RESULT resultid="1146" eventid="7" swimtime="00:00:38.01" lane="1" heatid="7008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="248" birthdate="2011-01-01" gender="F" lastname="Lekawska" firstname="Amelia" license="0">
              <RESULTS>
                <RESULT resultid="1147" eventid="5" swimtime="00:01:45.93" lane="2" heatid="5012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1148" eventid="7" swimtime="00:00:38.22" lane="4" heatid="7015" />
                <RESULT resultid="1149" eventid="19" swimtime="00:01:30.89" lane="1" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="249" birthdate="2010-01-01" gender="M" lastname="Malik" firstname="Adam" license="0">
              <RESULTS>
                <RESULT resultid="1150" eventid="8" status="DSQ" swimtime="00:00:30.97" lane="4" heatid="8020" comment="Der Sportler startete vor dem Startsignal" />
                <RESULT resultid="1151" eventid="14" swimtime="00:00:35.08" lane="1" heatid="14011" />
                <RESULT resultid="1152" eventid="18" swimtime="00:00:41.92" lane="1" heatid="18007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="250" birthdate="2013-01-01" gender="F" lastname="Mostowy" firstname="Maja" license="0">
              <RESULTS>
                <RESULT resultid="1153" eventid="3" swimtime="00:00:48.38" lane="2" heatid="3011" />
                <RESULT resultid="1154" eventid="7" swimtime="00:00:46.31" lane="2" heatid="7008" />
                <RESULT resultid="1155" eventid="17" swimtime="00:01:02.38" lane="3" heatid="17001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="251" birthdate="2013-01-01" gender="M" lastname="Nesterchuk" firstname="Mikolaj" license="0">
              <RESULTS>
                <RESULT resultid="1156" eventid="8" swimtime="00:00:33.29" lane="3" heatid="8005" />
                <RESULT resultid="1157" eventid="20" swimtime="00:01:16.79" lane="1" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="252" birthdate="2010-01-01" gender="M" lastname="Sieracki" firstname="Pawel" license="0">
              <RESULTS>
                <RESULT resultid="1158" eventid="8" swimtime="00:00:34.29" lane="2" heatid="8001" />
                <RESULT resultid="1159" eventid="14" status="DSQ" swimtime="00:00:46.70" lane="1" heatid="14001" comment="Der Sportler startete vor dem Startsignal" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="253" birthdate="2013-01-01" gender="F" lastname="Szurgot" firstname="Liliana" license="0">
              <RESULTS>
                <RESULT resultid="1160" eventid="7" swimtime="00:00:49.82" lane="1" heatid="7005" />
                <RESULT resultid="1161" eventid="17" swimtime="00:01:02.87" lane="2" heatid="17001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="254" birthdate="2012-01-01" gender="F" lastname="Szymkowicz" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="1162" eventid="3" status="DNS" swimtime="00:00:00.00" lane="1" heatid="3009" />
                <RESULT resultid="1163" eventid="7" status="DNS" swimtime="00:00:00.00" lane="3" heatid="7006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="255" birthdate="2011-01-01" gender="F" lastname="Szymkowicz" firstname="Maja" license="0">
              <RESULTS>
                <RESULT resultid="1164" eventid="3" swimtime="00:00:45.72" lane="2" heatid="3007" />
                <RESULT resultid="1165" eventid="7" swimtime="00:00:40.86" lane="4" heatid="7009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="256" birthdate="2012-01-01" gender="M" lastname="Tys" firstname="Wiktor" license="0">
              <RESULTS>
                <RESULT resultid="1166" eventid="8" swimtime="00:00:42.34" lane="2" heatid="8003" />
                <RESULT resultid="1167" eventid="18" swimtime="00:00:51.15" lane="3" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="257" birthdate="2011-01-01" gender="F" lastname="Wronkowska" firstname="Zofia" license="0">
              <RESULTS>
                <RESULT resultid="1168" eventid="3" swimtime="00:00:50.27" lane="4" heatid="3009" />
                <RESULT resultid="1169" eventid="7" swimtime="00:00:41.54" lane="2" heatid="7011" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Klub plavcu Melnickych" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="16" birthdate="2009-01-01" gender="F" lastname="Struplova" firstname="Ellen" license="0">
              <RESULTS>
                <RESULT resultid="65" eventid="31" swimtime="00:01:11.39" lane="1" heatid="31005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="66" eventid="33" swimtime="00:01:24.08" lane="2" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="67" eventid="43" swimtime="00:00:32.87" lane="3" heatid="43006" />
                <RESULT resultid="68" eventid="51" swimtime="00:02:33.26" lane="2" heatid="51004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="150" swimtime="00:01:54.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="17" birthdate="2009-01-01" gender="M" lastname="Zapp" firstname="Max" license="0">
              <RESULTS>
                <RESULT resultid="69" eventid="28" swimtime="00:00:35.74" lane="1" heatid="28006" />
                <RESULT resultid="70" eventid="32" swimtime="00:01:03.10" lane="2" heatid="32008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="71" eventid="38" swimtime="00:02:51.06" lane="2" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:22.26" />
                    <SPLIT distance="150" swimtime="00:02:06.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="72" eventid="44" swimtime="00:00:28.56" lane="2" heatid="44011" />
                <RESULT resultid="73" eventid="46" swimtime="00:01:18.26" lane="2" heatid="46003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="18" birthdate="2007-01-01" gender="F" lastname="Zloska" firstname="Karolina" license="0">
              <RESULTS>
                <RESULT resultid="74" eventid="31" swimtime="00:01:10.86" lane="2" heatid="31006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="75" eventid="33" swimtime="00:01:21.95" lane="4" heatid="33009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="76" eventid="41" swimtime="00:00:35.61" lane="1" heatid="41005" />
                <RESULT resultid="77" eventid="43" swimtime="00:00:32.84" lane="1" heatid="43009" />
                <RESULT resultid="78" eventid="53" swimtime="00:02:53.31" lane="3" heatid="53003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:21.61" />
                    <SPLIT distance="150" swimtime="00:02:15.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="19" birthdate="2006-01-01" gender="M" lastname="Zlosky" firstname="Adam" license="0">
              <RESULTS>
                <RESULT resultid="79" eventid="32" swimtime="00:00:56.31" lane="4" heatid="32010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="80" eventid="34" swimtime="00:01:07.03" lane="4" heatid="34007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="81" eventid="42" swimtime="00:00:28.02" lane="1" heatid="42007" />
                <RESULT resultid="82" eventid="44" swimtime="00:00:26.45" lane="2" heatid="44009" />
                <RESULT resultid="83" eventid="52" swimtime="00:02:04.62" lane="1" heatid="52005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="100" swimtime="00:01:00.36" />
                    <SPLIT distance="150" swimtime="00:01:32.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Neratovický plavecký klub" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="42" birthdate="2008-01-01" gender="M" lastname="Albert" firstname="Miroslav" license="56319000">
              <RESULTS>
                <RESULT resultid="153" eventid="26" swimtime="00:00:34.82" lane="3" heatid="26003" />
                <RESULT resultid="154" eventid="32" swimtime="00:01:07.20" lane="1" heatid="32004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="155" eventid="44" swimtime="00:00:30.17" lane="2" heatid="44003" />
                <RESULT resultid="156" eventid="48" swimtime="00:01:23.75" lane="3" heatid="48001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="157" eventid="52" swimtime="00:02:35.16" lane="2" heatid="52002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:13.27" />
                    <SPLIT distance="150" swimtime="00:01:56.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="43" birthdate="2011-01-01" gender="F" lastname="Brejchová" firstname="Eva" license="63441448">
              <RESULTS>
                <RESULT resultid="158" eventid="1" swimtime="00:01:41.32" lane="1" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="159" eventid="3" swimtime="00:00:41.48" lane="4" heatid="3022" />
                <RESULT resultid="160" eventid="7" swimtime="00:00:35.50" lane="2" heatid="7016" />
                <RESULT resultid="161" eventid="15" swimtime="00:01:29.24" lane="2" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="162" eventid="21" swimtime="00:03:13.16" lane="1" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                    <SPLIT distance="100" swimtime="00:01:33.95" />
                    <SPLIT distance="150" swimtime="00:02:30.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2008-01-01" gender="F" lastname="Broklová" firstname="Sofie" license="63440933">
              <RESULTS>
                <RESULT resultid="163" eventid="25" swimtime="00:00:40.61" lane="4" heatid="25003" />
                <RESULT resultid="164" eventid="31" swimtime="00:01:15.88" lane="3" heatid="31004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="165" eventid="33" swimtime="00:01:30.19" lane="4" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="166" eventid="41" swimtime="00:00:40.91" lane="1" heatid="41003" />
                <RESULT resultid="167" eventid="43" swimtime="00:00:33.59" lane="4" heatid="43006" />
                <RESULT resultid="168" eventid="47" swimtime="00:01:31.70" lane="4" heatid="47003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="45" birthdate="2004-01-01" gender="F" lastname="Dolanská" firstname="Johana" license="45991000">
              <RESULTS>
                <RESULT resultid="169" eventid="27" swimtime="00:00:38.14" lane="2" heatid="27009" />
                <RESULT resultid="170" eventid="31" swimtime="00:01:06.90" lane="4" heatid="31013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="171" eventid="37" swimtime="00:02:55.84" lane="4" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:02:09.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="172" eventid="41" swimtime="00:00:34.07" lane="4" heatid="41008" />
                <RESULT resultid="173" eventid="45" swimtime="00:01:23.04" lane="2" heatid="45007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="47" birthdate="2008-01-01" gender="M" lastname="Halász" firstname="Michal" license="56360000">
              <RESULTS>
                <RESULT resultid="179" eventid="30" swimtime="00:01:04.40" lane="1" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="180" eventid="32" swimtime="00:00:54.67" lane="3" heatid="32009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="181" eventid="42" swimtime="00:00:27.79" lane="1" heatid="42010" />
                <RESULT resultid="182" eventid="44" swimtime="00:00:24.60" lane="3" heatid="44012" />
                <RESULT resultid="183" eventid="52" swimtime="00:02:07.41" lane="4" heatid="52005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="100" swimtime="00:01:01.38" />
                    <SPLIT distance="150" swimtime="00:01:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2082" eventid="65" swimtime="00:00:26.72" lane="4" heatid="65001" />
                <RESULT resultid="2096" eventid="69" swimtime="00:00:24.46" lane="2" heatid="69001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="48" birthdate="2008-01-01" gender="F" lastname="Hnátková" firstname="Johana" license="51814000">
              <RESULTS>
                <RESULT resultid="184" eventid="25" swimtime="00:00:35.64" lane="1" heatid="25006" />
                <RESULT resultid="185" eventid="31" swimtime="00:01:07.65" lane="1" heatid="31008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="186" eventid="35" swimtime="00:02:44.87" lane="2" heatid="35002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:20.08" />
                    <SPLIT distance="150" swimtime="00:02:04.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="187" eventid="43" swimtime="00:00:30.57" lane="3" heatid="43010" />
                <RESULT resultid="188" eventid="51" swimtime="00:02:25.84" lane="1" heatid="51005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:09.51" />
                    <SPLIT distance="150" swimtime="00:01:49.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="49" birthdate="2005-01-01" gender="F" lastname="Hrdinová" firstname="Natálie" license="37833000">
              <RESULTS>
                <RESULT resultid="189" eventid="29" swimtime="00:01:17.71" lane="3" heatid="29006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="190" eventid="37" swimtime="00:03:02.28" lane="1" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                    <SPLIT distance="100" swimtime="00:01:27.00" />
                    <SPLIT distance="150" swimtime="00:02:14.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="191" eventid="45" swimtime="00:01:24.88" lane="1" heatid="45006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="192" eventid="49" swimtime="00:02:46.59" lane="1" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:18.71" />
                    <SPLIT distance="150" swimtime="00:02:02.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="50" birthdate="2007-01-01" gender="F" lastname="Lipenská" firstname="Klára" license="40345000">
              <RESULTS>
                <RESULT resultid="193" eventid="29" swimtime="00:01:11.21" lane="3" heatid="29005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="194" eventid="31" swimtime="00:01:02.00" lane="2" heatid="31011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="195" eventid="41" swimtime="00:00:31.36" lane="4" heatid="41012" />
                <RESULT resultid="196" eventid="43" swimtime="00:00:28.04" lane="3" heatid="43015" />
                <RESULT resultid="197" eventid="51" swimtime="00:02:16.68" lane="3" heatid="51005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:05.54" />
                    <SPLIT distance="150" swimtime="00:01:41.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2072" eventid="63" swimtime="00:00:31.01" lane="3" heatid="63001" />
                <RESULT resultid="2088" eventid="67" swimtime="00:00:27.89" lane="3" heatid="67001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="51" birthdate="2008-01-01" gender="M" lastname="Novák" firstname="Matyás" license="51406000">
              <RESULTS>
                <RESULT resultid="198" eventid="28" swimtime="00:00:35.92" lane="2" heatid="28002" />
                <RESULT resultid="199" eventid="32" swimtime="00:01:04.88" lane="2" heatid="32004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="200" eventid="44" swimtime="00:00:30.26" lane="4" heatid="44004" />
                <RESULT resultid="201" eventid="46" swimtime="00:01:20.29" lane="4" heatid="46004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="202" eventid="54" swimtime="00:02:42.33" lane="4" heatid="54002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:16.79" />
                    <SPLIT distance="150" swimtime="00:02:02.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="52" birthdate="2007-01-01" gender="F" lastname="Salajková" firstname="Mariana" license="45351000">
              <RESULTS>
                <RESULT resultid="203" eventid="27" swimtime="00:00:40.60" lane="1" heatid="27004" />
                <RESULT resultid="204" eventid="31" swimtime="00:01:13.53" lane="4" heatid="31005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="205" eventid="37" swimtime="00:03:15.43" lane="1" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:32.00" />
                    <SPLIT distance="150" swimtime="00:02:24.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="206" eventid="43" swimtime="00:00:33.41" lane="1" heatid="43006" />
                <RESULT resultid="207" eventid="45" swimtime="00:01:31.15" lane="3" heatid="45002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="53" birthdate="2010-01-01" gender="M" lastname="Tichý" firstname="Simon" license="63440889">
              <RESULTS>
                <RESULT resultid="208" eventid="2" status="DNS" swimtime="00:00:00.00" lane="2" heatid="2004" />
                <RESULT resultid="209" eventid="4" status="DNS" swimtime="00:00:00.00" lane="4" heatid="4015" />
                <RESULT resultid="210" eventid="14" status="DNS" swimtime="00:00:00.00" lane="2" heatid="14006" />
                <RESULT resultid="211" eventid="18" status="DNS" swimtime="00:00:00.00" lane="4" heatid="18013" />
                <RESULT resultid="212" eventid="20" status="DNS" swimtime="00:00:00.00" lane="2" heatid="20010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="54" birthdate="2014-01-01" gender="M" lastname="Tvrdík" firstname="Matteo" license="63456334">
              <RESULTS>
                <RESULT resultid="213" eventid="6" swimtime="00:02:01.74" lane="3" heatid="6006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="214" eventid="8" swimtime="00:00:42.94" lane="2" heatid="8004" />
                <RESULT resultid="215" eventid="10" swimtime="00:02:01.37" lane="2" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="216" eventid="18" status="DSQ" swimtime="00:00:54.09" lane="1" heatid="18009" comment="Der Sportler startete vor dem Startsignal" />
                <RESULT resultid="217" eventid="20" swimtime="00:01:41.64" lane="3" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="55" birthdate="2008-01-01" gender="M" lastname="Valko" firstname="Jakub" license="45172000">
              <RESULTS>
                <RESULT resultid="218" eventid="26" swimtime="00:00:32.28" lane="3" heatid="26004" />
                <RESULT resultid="219" eventid="28" swimtime="00:00:35.91" lane="3" heatid="28003" />
                <RESULT resultid="220" eventid="34" swimtime="00:01:10.97" lane="3" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="221" eventid="44" swimtime="00:00:27.13" lane="3" heatid="44006" />
                <RESULT resultid="222" eventid="52" swimtime="00:02:13.62" lane="4" heatid="52004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="150" swimtime="00:01:36.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="56" birthdate="2008-01-01" gender="M" lastname="Zaludek" firstname="Martin" license="43542000">
              <RESULTS>
                <RESULT resultid="223" eventid="28" swimtime="00:00:33.83" lane="3" heatid="28004" />
                <RESULT resultid="224" eventid="32" swimtime="00:01:00.63" lane="3" heatid="32006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="225" eventid="42" swimtime="00:00:30.42" lane="3" heatid="42004" />
                <RESULT resultid="226" eventid="44" swimtime="00:00:27.26" lane="1" heatid="44007" />
                <RESULT resultid="227" eventid="52" swimtime="00:02:18.41" lane="3" heatid="52004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:04.65" />
                    <SPLIT distance="150" swimtime="00:01:42.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1946" eventid="40" swimtime="00:01:49.22" lane="1" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.56" />
                    <SPLIT distance="100" swimtime="00:00:51.53" />
                    <SPLIT distance="150" swimtime="00:01:20.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47" number="1" />
                    <RELAYPOSITION athleteid="55" number="2" />
                    <RELAYPOSITION athleteid="42" number="3" />
                    <RELAYPOSITION athleteid="51" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1947" eventid="72" swimtime="00:02:01.09" lane="2" heatid="72001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:01:05.83" />
                    <SPLIT distance="150" swimtime="00:01:33.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="55" number="1" />
                    <RELAYPOSITION athleteid="56" number="2" />
                    <RELAYPOSITION athleteid="47" number="3" />
                    <RELAYPOSITION athleteid="51" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1948" eventid="39" swimtime="00:02:07.09" lane="2" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:01.23" />
                    <SPLIT distance="150" swimtime="00:01:34.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48" number="1" />
                    <RELAYPOSITION athleteid="49" number="2" />
                    <RELAYPOSITION athleteid="44" number="3" />
                    <RELAYPOSITION athleteid="52" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1949" eventid="71" swimtime="00:02:15.50" lane="2" heatid="71001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:13.18" />
                    <SPLIT distance="150" swimtime="00:01:46.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48" number="1" />
                    <RELAYPOSITION athleteid="45" number="2" />
                    <RELAYPOSITION athleteid="49" number="3" />
                    <RELAYPOSITION athleteid="50" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Plavecký klub Litvínov" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="58" birthdate="2013-01-01" gender="M" lastname="Geier" firstname="Sebastian" license="0">
              <RESULTS>
                <RESULT resultid="232" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="233" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="234" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="235" eventid="20" status="WDR" swimtime="00:00:00.00" lane="0" heatid="20000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="59" birthdate="2014-01-01" gender="M" lastname="Gergel" firstname="Adam" license="0">
              <RESULTS>
                <RESULT resultid="236" eventid="4" swimtime="00:00:49.22" lane="3" heatid="4002" />
                <RESULT resultid="237" eventid="8" swimtime="00:00:46.22" lane="3" heatid="8003" />
                <RESULT resultid="238" eventid="16" swimtime="00:01:53.38" lane="2" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="239" eventid="20" swimtime="00:01:51.06" lane="3" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="60" birthdate="2012-01-01" gender="F" lastname="Kejrová" firstname="Lucie" license="0">
              <RESULTS>
                <RESULT resultid="240" eventid="1" swimtime="00:01:39.80" lane="2" heatid="1001">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:44.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="241" eventid="9" swimtime="00:01:36.22" lane="1" heatid="9008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="242" eventid="13" swimtime="00:00:43.63" lane="1" heatid="13005" />
                <RESULT resultid="243" eventid="15" swimtime="00:01:33.14" lane="1" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="61" birthdate="2012-01-01" gender="F" lastname="Kejrová" firstname="Markéta" license="0">
              <RESULTS>
                <RESULT resultid="244" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="245" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="246" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="247" eventid="19" status="WDR" swimtime="00:00:00.00" lane="0" heatid="19000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="62" birthdate="2013-01-01" gender="M" lastname="Kovarik" firstname="Jakub" license="0">
              <RESULTS>
                <RESULT resultid="248" eventid="6" swimtime="00:01:36.64" lane="3" heatid="6007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="249" eventid="10" swimtime="00:01:27.61" lane="1" heatid="10008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="250" eventid="14" swimtime="00:00:41.96" lane="3" heatid="14005" />
                <RESULT resultid="251" eventid="18" swimtime="00:00:43.85" lane="2" heatid="18010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="63" birthdate="2013-01-01" gender="F" lastname="Langhammerová" firstname="Ella" license="0">
              <RESULTS>
                <RESULT resultid="252" eventid="3" status="WDR" swimtime="00:00:00.00" lane="0" heatid="3000" />
                <RESULT resultid="253" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="254" eventid="15" status="WDR" swimtime="00:00:00.00" lane="0" heatid="15000" />
                <RESULT resultid="255" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="64" birthdate="2008-01-01" gender="F" lastname="Lisková" firstname="Julie" license="0">
              <RESULTS>
                <RESULT resultid="256" eventid="27" swimtime="00:00:38.94" lane="2" heatid="27004" />
                <RESULT resultid="257" eventid="37" swimtime="00:03:05.53" lane="2" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:29.65" />
                    <SPLIT distance="150" swimtime="00:02:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="258" eventid="45" swimtime="00:01:26.05" lane="2" heatid="45002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="259" eventid="53" swimtime="00:02:55.66" lane="2" heatid="53002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:25.49" />
                    <SPLIT distance="150" swimtime="00:02:14.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2056" eventid="59" swimtime="00:00:38.66" lane="4" heatid="59001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="66" birthdate="2013-01-01" gender="F" lastname="Pechová" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="262" eventid="3" swimtime="00:00:39.80" lane="1" heatid="3020" />
                <RESULT resultid="263" eventid="7" swimtime="00:00:35.45" lane="1" heatid="7021" />
                <RESULT resultid="264" eventid="15" swimtime="00:01:29.88" lane="3" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="265" eventid="19" swimtime="00:01:23.60" lane="3" heatid="19014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="67" birthdate="2008-01-01" gender="F" lastname="Prantová" firstname="Laura" license="0">
              <RESULTS>
                <RESULT resultid="266" eventid="25" swimtime="00:00:32.55" lane="3" heatid="25011" />
                <RESULT resultid="267" eventid="29" swimtime="00:01:13.38" lane="4" heatid="29005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="268" eventid="41" swimtime="00:00:31.63" lane="2" heatid="41009" />
                <RESULT resultid="269" eventid="43" swimtime="00:00:29.79" lane="4" heatid="43012" />
                <RESULT resultid="2039" eventid="55" swimtime="00:00:32.81" lane="1" heatid="55001" />
                <RESULT resultid="2073" eventid="63" swimtime="00:00:31.34" lane="1" heatid="63001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="68" birthdate="2011-01-01" gender="F" lastname="Praská" firstname="Adéla" license="0">
              <RESULTS>
                <RESULT resultid="270" eventid="5" swimtime="00:01:35.94" lane="1" heatid="5007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="271" eventid="7" swimtime="00:00:33.91" lane="4" heatid="7018" />
                <RESULT resultid="272" eventid="15" swimtime="00:01:31.65" lane="3" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="273" eventid="21" swimtime="00:03:11.39" lane="2" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                    <SPLIT distance="100" swimtime="00:01:37.98" />
                    <SPLIT distance="150" swimtime="00:02:31.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="69" birthdate="2012-01-01" gender="F" lastname="Raciková" firstname="Hana" license="0">
              <RESULTS>
                <RESULT resultid="274" eventid="5" swimtime="00:01:35.19" lane="4" heatid="5011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="275" eventid="7" swimtime="00:00:34.75" lane="1" heatid="7017" />
                <RESULT resultid="276" eventid="15" swimtime="00:01:24.82" lane="3" heatid="15013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="277" eventid="21" swimtime="00:03:02.15" lane="3" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:27.32" />
                    <SPLIT distance="150" swimtime="00:02:19.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="70" birthdate="2008-01-01" gender="M" lastname="Rous" firstname="David" license="0">
              <RESULTS>
                <RESULT resultid="278" eventid="26" swimtime="00:00:29.99" lane="1" heatid="26009" />
                <RESULT resultid="279" eventid="32" swimtime="00:00:57.96" lane="4" heatid="32009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="280" eventid="42" swimtime="00:00:28.52" lane="4" heatid="42006" />
                <RESULT resultid="281" eventid="48" swimtime="00:01:06.28" lane="1" heatid="48004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="71" birthdate="2012-01-01" gender="F" lastname="Rovná" firstname="Julie" license="0">
              <RESULTS>
                <RESULT resultid="282" eventid="5" swimtime="00:01:49.31" lane="1" heatid="5005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="283" eventid="7" swimtime="00:00:41.53" lane="1" heatid="7011" />
                <RESULT resultid="284" eventid="13" swimtime="00:00:53.14" lane="3" heatid="13002" />
                <RESULT resultid="285" eventid="15" swimtime="00:01:44.78" lane="2" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="72" birthdate="2008-01-01" gender="M" lastname="Stafa" firstname="Pavel" license="0">
              <RESULTS>
                <RESULT resultid="286" eventid="26" status="DNS" swimtime="00:00:00.00" lane="4" heatid="26004" />
                <RESULT resultid="287" eventid="32" status="DNS" swimtime="00:00:00.00" lane="1" heatid="32005" />
                <RESULT resultid="288" eventid="44" status="DNS" swimtime="00:00:00.00" lane="3" heatid="44005" />
                <RESULT resultid="289" eventid="48" status="DNS" swimtime="00:00:00.00" lane="1" heatid="48002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="73" birthdate="2011-01-01" gender="F" lastname="Struharonská" firstname="Alica" license="0">
              <RESULTS>
                <RESULT resultid="290" eventid="1" swimtime="00:01:28.44" lane="3" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="291" eventid="7" swimtime="00:00:32.90" lane="1" heatid="7018" />
                <RESULT resultid="292" eventid="15" swimtime="00:01:24.50" lane="4" heatid="15014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="293" eventid="21" swimtime="00:03:07.48" lane="2" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                    <SPLIT distance="100" swimtime="00:01:29.09" />
                    <SPLIT distance="150" swimtime="00:02:25.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="74" birthdate="2013-01-01" gender="F" lastname="Ulrichová" firstname="Eliska" license="0">
              <RESULTS>
                <RESULT resultid="294" eventid="5" status="WDR" swimtime="00:00:00.00" lane="0" heatid="5000" />
                <RESULT resultid="295" eventid="9" status="WDR" swimtime="00:00:00.00" lane="0" heatid="9000" />
                <RESULT resultid="296" eventid="13" status="WDR" swimtime="00:00:00.00" lane="0" heatid="13000" />
                <RESULT resultid="297" eventid="17" status="WDR" swimtime="00:00:00.00" lane="0" heatid="17000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="75" birthdate="2013-01-01" gender="M" lastname="Vojtuloviè" firstname="Filip" license="0">
              <RESULTS>
                <RESULT resultid="298" eventid="2" swimtime="00:01:44.26" lane="2" heatid="2001">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:48.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="299" eventid="10" swimtime="00:01:36.46" lane="4" heatid="10008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="300" eventid="14" swimtime="00:00:42.03" lane="4" heatid="14008" />
                <RESULT resultid="301" eventid="20" swimtime="00:01:25.15" lane="1" heatid="20009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="76" birthdate="2015-01-01" gender="F" lastname="Vojtulovièová" firstname="Ema" license="0">
              <RESULTS>
                <RESULT resultid="302" eventid="3" swimtime="00:00:54.66" lane="3" heatid="3002" />
                <RESULT resultid="303" eventid="7" swimtime="00:00:59.26" lane="2" heatid="7001" />
                <RESULT resultid="304" eventid="17" swimtime="00:01:05.55" lane="4" heatid="17002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="77" birthdate="2012-01-01" gender="M" lastname="Zicha" firstname="Pavel" license="0">
              <RESULTS>
                <RESULT resultid="305" eventid="2" swimtime="00:01:22.07" lane="3" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="306" eventid="6" swimtime="00:01:30.86" lane="1" heatid="6008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="307" eventid="14" swimtime="00:00:34.96" lane="1" heatid="14009" />
                <RESULT resultid="308" eventid="20" swimtime="00:01:09.08" lane="1" heatid="20014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="260" eventid="11" swimtime="00:02:10.93" lane="3" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:40.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="73" number="1" />
                    <RELAYPOSITION athleteid="69" number="2" />
                    <RELAYPOSITION athleteid="62" number="3" />
                    <RELAYPOSITION athleteid="77" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="261" eventid="23" swimtime="00:02:30.42" lane="3" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:01:56.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="69" number="1" />
                    <RELAYPOSITION athleteid="62" number="2" />
                    <RELAYPOSITION athleteid="77" number="3" />
                    <RELAYPOSITION athleteid="73" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Plavecky klub Most" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="106" birthdate="2010-01-01" gender="M" lastname="Augustín" firstname="Tomás" license="0">
              <RESULTS>
                <RESULT resultid="440" eventid="4" swimtime="00:00:33.41" lane="2" heatid="4015" />
                <RESULT resultid="441" eventid="8" swimtime="00:00:28.65" lane="3" heatid="8020" />
                <RESULT resultid="442" eventid="10" swimtime="00:01:14.85" lane="3" heatid="10011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="443" eventid="14" swimtime="00:00:31.78" lane="3" heatid="14011" />
                <RESULT resultid="444" eventid="20" swimtime="00:01:04.27" lane="3" heatid="20016">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="2013-01-01" gender="F" lastname="Behrová" firstname="Nicol" license="0">
              <RESULTS>
                <RESULT resultid="445" eventid="3" swimtime="00:00:52.06" lane="4" heatid="3008" />
                <RESULT resultid="446" eventid="7" swimtime="00:00:47.22" lane="4" heatid="7007" />
                <RESULT resultid="447" eventid="9" status="DNS" swimtime="00:00:00.00" lane="4" heatid="9004" />
                <RESULT resultid="448" eventid="15" swimtime="00:01:50.56" lane="1" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="449" eventid="19" swimtime="00:01:44.58" lane="3" heatid="19004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2013-01-01" gender="F" lastname="Boudníková" firstname="Lucie" license="0">
              <RESULTS>
                <RESULT resultid="450" eventid="5" status="DNS" swimtime="00:00:00.00" lane="3" heatid="5010" />
                <RESULT resultid="451" eventid="7" status="DNS" swimtime="00:00:00.00" lane="3" heatid="7021" />
                <RESULT resultid="452" eventid="9" status="DNS" swimtime="00:00:00.00" lane="2" heatid="9013" />
                <RESULT resultid="453" eventid="17" status="DNS" swimtime="00:00:00.00" lane="3" heatid="17012" />
                <RESULT resultid="454" eventid="21" status="DNS" swimtime="00:00:00.00" lane="1" heatid="21004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="2008-01-01" gender="M" lastname="Brázda" firstname="Ondrej" license="0">
              <RESULTS>
                <RESULT resultid="455" eventid="28" swimtime="00:00:41.66" lane="2" heatid="28001" />
                <RESULT resultid="456" eventid="34" swimtime="00:01:17.95" lane="4" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="457" eventid="42" swimtime="00:00:31.70" lane="2" heatid="42004" />
                <RESULT resultid="458" eventid="44" swimtime="00:00:30.12" lane="4" heatid="44006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110" birthdate="2004-01-01" gender="F" lastname="Cervinková" firstname="Emma" license="0">
              <RESULTS>
                <RESULT resultid="459" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
                <RESULT resultid="460" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="461" eventid="31" status="WDR" swimtime="00:00:00.00" lane="0" heatid="31000" />
                <RESULT resultid="462" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
                <RESULT resultid="463" eventid="45" status="WDR" swimtime="00:00:00.00" lane="0" heatid="45000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111" birthdate="2009-01-01" gender="F" lastname="Dunková" firstname="Helena" license="0">
              <RESULTS>
                <RESULT resultid="464" eventid="25" swimtime="00:00:38.43" lane="4" heatid="25005" />
                <RESULT resultid="465" eventid="27" swimtime="00:00:41.93" lane="4" heatid="27003" />
                <RESULT resultid="466" eventid="33" swimtime="00:01:22.25" lane="4" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="467" eventid="41" swimtime="00:00:35.28" lane="4" heatid="41006" />
                <RESULT resultid="468" eventid="43" swimtime="00:00:33.07" lane="3" heatid="43007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="112" birthdate="2012-01-01" gender="F" lastname="Maksymiv" firstname="Lilija" license="0">
              <RESULTS>
                <RESULT resultid="469" eventid="5" swimtime="00:01:51.67" lane="4" heatid="5004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="470" eventid="7" swimtime="00:00:42.13" lane="3" heatid="7011" />
                <RESULT resultid="471" eventid="9" swimtime="00:01:49.96" lane="4" heatid="9006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="472" eventid="19" swimtime="00:01:35.22" lane="2" heatid="19006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113" birthdate="2009-01-01" gender="M" lastname="Najmon" firstname="Tomás" license="0">
              <RESULTS>
                <RESULT resultid="473" eventid="28" swimtime="00:00:36.55" lane="4" heatid="28006" />
                <RESULT resultid="474" eventid="32" swimtime="00:01:06.89" lane="2" heatid="32003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="475" eventid="38" swimtime="00:03:00.21" lane="1" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:02:12.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="476" eventid="44" swimtime="00:00:29.98" lane="1" heatid="44011" />
                <RESULT resultid="477" eventid="46" swimtime="00:01:20.47" lane="4" heatid="46003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="114" birthdate="2011-01-01" gender="F" lastname="Rejmanová" firstname="Barbora" license="0">
              <RESULTS>
                <RESULT resultid="478" eventid="3" swimtime="00:00:43.72" lane="1" heatid="3015" />
                <RESULT resultid="479" eventid="7" swimtime="00:00:35.81" lane="2" heatid="7015" />
                <RESULT resultid="480" eventid="9" swimtime="00:01:35.50" lane="3" heatid="9008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="481" eventid="15" swimtime="00:01:36.78" lane="1" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="482" eventid="19" swimtime="00:01:21.69" lane="3" heatid="19009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="115" birthdate="2014-01-01" gender="M" lastname="Rychlý" firstname="Jan" license="0">
              <RESULTS>
                <RESULT resultid="483" eventid="4" swimtime="00:00:37.82" lane="2" heatid="4011" />
                <RESULT resultid="484" eventid="8" swimtime="00:00:32.57" lane="2" heatid="8016" />
                <RESULT resultid="485" eventid="14" swimtime="00:00:37.38" lane="2" heatid="14007" />
                <RESULT resultid="486" eventid="20" swimtime="00:01:14.15" lane="2" heatid="20012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="116" birthdate="2014-01-01" gender="M" lastname="Vacek" firstname="Jáchym" license="0">
              <RESULTS>
                <RESULT resultid="487" eventid="4" swimtime="00:00:42.00" lane="3" heatid="4011" />
                <RESULT resultid="488" eventid="8" swimtime="00:00:35.03" lane="1" heatid="8016" />
                <RESULT resultid="489" eventid="16" status="DSQ" swimtime="00:01:30.81" lane="3" heatid="16005" comment="Der Sportler hat bei der dritten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="490" eventid="18" status="DSQ" swimtime="00:00:50.27" lane="2" heatid="18009" comment="Nach der Wende  hat der Sportler zwei Delphinbeinschläge ausgeführt." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="117" birthdate="2014-01-01" gender="M" lastname="Valenta" firstname="Krystof" license="0">
              <RESULTS>
                <RESULT resultid="491" eventid="4" swimtime="00:00:45.45" lane="4" heatid="4006" />
                <RESULT resultid="492" eventid="8" swimtime="00:00:39.73" lane="1" heatid="8006" />
                <RESULT resultid="493" eventid="14" status="DSQ" swimtime="00:00:50.18" lane="4" heatid="14007" comment="Der Sportler führte mit den Beinen auf der Schwimmstrecke wechselseitig Bewegungen aus." />
                <RESULT resultid="494" eventid="20" swimtime="00:01:28.11" lane="1" heatid="20012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Aqua Köln" nation="GER" region="17" code="6449">
          <ATHLETES>
            <ATHLETE athleteid="20" birthdate="1993-01-01" gender="M" lastname="Felsner" firstname="Stefan" license="147637">
              <RESULTS>
                <RESULT resultid="84" eventid="26" status="DNS" swimtime="00:00:00.00" lane="4" heatid="26011" />
                <RESULT resultid="85" eventid="30" swimtime="00:00:55.84" lane="2" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="86" eventid="42" swimtime="00:00:25.32" lane="3" heatid="42012" />
                <RESULT resultid="87" eventid="44" swimtime="00:00:23.74" lane="3" heatid="44014" />
                <RESULT resultid="2084" eventid="66" swimtime="00:00:25.28" lane="3" heatid="66001" />
                <RESULT resultid="2101" eventid="70" swimtime="00:00:23.60" lane="3" heatid="70001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Chemnitz von 1892" nation="GER" region="12" code="3353">
          <ATHLETES>
            <ATHLETE athleteid="101" birthdate="2011-01-01" gender="F" lastname="Franke" firstname="Loreley" license="447682">
              <RESULTS>
                <RESULT resultid="413" eventid="3" swimtime="00:00:35.28" lane="3" heatid="3022" />
                <RESULT resultid="414" eventid="7" swimtime="00:00:31.39" lane="1" heatid="7023" />
                <RESULT resultid="415" eventid="15" swimtime="00:01:19.13" lane="3" heatid="15014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="416" eventid="19" swimtime="00:01:08.57" lane="3" heatid="19016">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="417" eventid="35" swimtime="00:02:47.69" lane="1" heatid="35002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:20.17" />
                    <SPLIT distance="150" swimtime="00:02:04.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="418" eventid="51" swimtime="00:02:36.81" lane="1" heatid="51004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                    <SPLIT distance="150" swimtime="00:01:57.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102" birthdate="2005-01-01" gender="F" lastname="Furka" firstname="Vanessa" license="351356">
              <RESULTS>
                <RESULT resultid="419" eventid="25" swimtime="00:00:30.18" lane="2" heatid="25012" />
                <RESULT resultid="420" eventid="31" swimtime="00:00:59.94" lane="2" heatid="31012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="421" eventid="41" swimtime="00:00:29.43" lane="3" heatid="41013" />
                <RESULT resultid="422" eventid="43" swimtime="00:00:27.69" lane="3" heatid="43016" />
                <RESULT resultid="423" eventid="53" swimtime="00:02:30.76" lane="1" heatid="53005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:56.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2042" eventid="56" swimtime="00:00:30.58" lane="3" heatid="56001" />
                <RESULT resultid="2078" eventid="64" swimtime="00:00:28.95" lane="4" heatid="64001" />
                <RESULT resultid="2094" eventid="68" swimtime="00:00:27.58" lane="4" heatid="68001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="103" birthdate="2012-01-01" gender="M" lastname="Gehre" firstname="Matti" license="437418">
              <RESULTS>
                <RESULT resultid="424" eventid="4" swimtime="00:00:38.44" lane="4" heatid="4013" />
                <RESULT resultid="425" eventid="8" swimtime="00:00:31.69" lane="3" heatid="8018" />
                <RESULT resultid="426" eventid="16" swimtime="00:01:24.14" lane="1" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="427" eventid="20" swimtime="00:01:10.72" lane="2" heatid="20014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="428" eventid="36" swimtime="00:02:59.40" lane="1" heatid="36001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                    <SPLIT distance="100" swimtime="00:01:29.65" />
                    <SPLIT distance="150" swimtime="00:02:16.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="429" eventid="52" swimtime="00:02:36.10" lane="1" heatid="52003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="150" swimtime="00:01:56.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="104" birthdate="2013-01-01" gender="M" lastname="Goebel" firstname="Ferdinand" license="444239">
              <RESULTS>
                <RESULT resultid="430" eventid="6" swimtime="00:01:32.48" lane="2" heatid="6007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="431" eventid="8" swimtime="00:00:32.99" lane="4" heatid="8011" />
                <RESULT resultid="432" eventid="14" swimtime="00:00:37.30" lane="3" heatid="14006" />
                <RESULT resultid="433" eventid="20" swimtime="00:01:13.72" lane="4" heatid="20013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="434" eventid="38" status="DNS" swimtime="00:00:00.00" lane="3" heatid="38001" />
                <RESULT resultid="435" eventid="52" status="DNS" swimtime="00:00:00.00" lane="2" heatid="52001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105" birthdate="2005-01-01" gender="F" lastname="Prochaska" firstname="Susanna" license="325221">
              <RESULTS>
                <RESULT resultid="436" eventid="25" status="WDR" swimtime="00:00:00.00" lane="0" heatid="25000" />
                <RESULT resultid="437" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="438" eventid="33" status="WDR" swimtime="00:00:00.00" lane="0" heatid="33000" />
                <RESULT resultid="439" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Eintracht Berlin e.V." nation="GER" region="3" code="5673">
          <ATHLETES>
            <ATHLETE athleteid="82" birthdate="2012-01-01" gender="F" lastname="Baumert" firstname="Lisa" license="463365">
              <RESULTS>
                <RESULT resultid="314" eventid="3" status="DNS" swimtime="00:00:00.00" lane="2" heatid="3009" />
                <RESULT resultid="315" eventid="7" status="DNS" swimtime="00:00:00.00" lane="3" heatid="7007" />
                <RESULT resultid="316" eventid="9" status="DNS" swimtime="00:00:00.00" lane="4" heatid="9005" />
                <RESULT resultid="317" eventid="17" status="DNS" swimtime="00:00:00.00" lane="1" heatid="17005" />
                <RESULT resultid="318" eventid="19" status="DNS" swimtime="00:00:00.00" lane="4" heatid="19003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="83" birthdate="2011-01-01" gender="F" lastname="Baumert" firstname="Marie" license="450130">
              <RESULTS>
                <RESULT resultid="319" eventid="3" swimtime="00:00:46.70" lane="3" heatid="3010" />
                <RESULT resultid="320" eventid="5" swimtime="00:01:47.18" lane="4" heatid="5003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="321" eventid="9" swimtime="00:01:41.60" lane="1" heatid="9006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="322" eventid="19" swimtime="00:01:36.91" lane="4" heatid="19004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="323" eventid="37" status="DNS" swimtime="00:00:00.00" lane="1" heatid="37001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="84" birthdate="2009-01-01" gender="F" lastname="Cappelli" firstname="Emma" license="386111">
              <RESULTS>
                <RESULT resultid="324" eventid="31" swimtime="00:01:08.04" lane="2" heatid="31004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="325" eventid="33" swimtime="00:01:18.89" lane="1" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="326" eventid="41" swimtime="00:00:33.50" lane="3" heatid="41006" />
                <RESULT resultid="327" eventid="43" swimtime="00:00:30.43" lane="3" heatid="43011" />
                <RESULT resultid="328" eventid="51" swimtime="00:02:42.66" lane="2" heatid="51003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:02:05.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="85" birthdate="2005-01-01" gender="M" lastname="Deister" firstname="Marvin" license="327479">
              <RESULTS>
                <RESULT resultid="329" eventid="26" status="DNS" swimtime="00:00:00.00" lane="2" heatid="26006" />
                <RESULT resultid="330" eventid="28" status="WDR" swimtime="00:00:00.00" lane="0" heatid="28000" />
                <RESULT resultid="331" eventid="32" status="DNS" swimtime="00:00:00.00" lane="2" heatid="32006" />
                <RESULT resultid="332" eventid="42" status="DNS" swimtime="00:00:00.00" lane="1" heatid="42011" />
                <RESULT resultid="333" eventid="44" status="DNS" swimtime="00:00:00.00" lane="4" heatid="44013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="86" birthdate="2010-01-01" gender="F" lastname="Dorn" firstname="Anne" license="435621">
              <RESULTS>
                <RESULT resultid="334" eventid="27" swimtime="00:00:41.18" lane="3" heatid="27005" />
                <RESULT resultid="335" eventid="31" swimtime="00:01:19.31" lane="1" heatid="31001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="336" eventid="41" swimtime="00:00:43.68" lane="2" heatid="41001" />
                <RESULT resultid="337" eventid="43" swimtime="00:00:34.77" lane="1" heatid="43005" />
                <RESULT resultid="338" eventid="51" swimtime="00:03:06.48" lane="2" heatid="51002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:29.10" />
                    <SPLIT distance="150" swimtime="00:02:19.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="87" birthdate="2011-01-01" gender="M" lastname="Feige" firstname="Bennet" license="441662">
              <RESULTS>
                <RESULT resultid="339" eventid="4" swimtime="00:00:45.08" lane="3" heatid="4005" />
                <RESULT resultid="340" eventid="8" swimtime="00:00:36.73" lane="3" heatid="8009" />
                <RESULT resultid="341" eventid="10" swimtime="00:01:38.77" lane="4" heatid="10010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="342" eventid="14" swimtime="00:00:48.04" lane="3" heatid="14003" />
                <RESULT resultid="343" eventid="20" swimtime="00:01:27.68" lane="4" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="88" birthdate="2007-01-01" gender="M" lastname="Hahn" firstname="Artur" license="386117">
              <RESULTS>
                <RESULT resultid="344" eventid="26" swimtime="00:00:36.35" lane="3" heatid="26002" />
                <RESULT resultid="345" eventid="32" swimtime="00:01:09.28" lane="2" heatid="32002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="346" eventid="42" swimtime="00:00:34.47" lane="3" heatid="42001" />
                <RESULT resultid="347" eventid="44" swimtime="00:00:30.44" lane="2" heatid="44004" />
                <RESULT resultid="348" eventid="48" swimtime="00:01:22.72" lane="2" heatid="48001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="89" birthdate="2010-01-01" gender="F" lastname="Hinze" firstname="Frieda Luise" license="425043">
              <RESULTS>
                <RESULT resultid="349" eventid="27" status="DSQ" swimtime="00:00:45.22" lane="4" heatid="27005" comment="Nach dem Start hat der Sportler zwei Tauchzüge ausgeführt." />
                <RESULT resultid="350" eventid="31" swimtime="00:01:28.87" lane="3" heatid="31001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="351" eventid="33" swimtime="00:01:36.11" lane="3" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="352" eventid="41" swimtime="00:00:41.42" lane="1" heatid="41002" />
                <RESULT resultid="353" eventid="43" swimtime="00:00:39.07" lane="2" heatid="43001" />
                <RESULT resultid="354" eventid="53" swimtime="00:03:34.75" lane="1" heatid="53002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                    <SPLIT distance="100" swimtime="00:01:39.66" />
                    <SPLIT distance="150" swimtime="00:02:41.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="90" birthdate="2014-01-01" gender="F" lastname="Kallinich" firstname="Marie" license="467500">
              <RESULTS>
                <RESULT resultid="355" eventid="3" swimtime="00:00:44.19" lane="1" heatid="3010" />
                <RESULT resultid="356" eventid="7" swimtime="00:00:41.72" lane="3" heatid="7008" />
                <RESULT resultid="357" eventid="9" swimtime="00:01:44.45" lane="1" heatid="9004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="358" eventid="15" swimtime="00:01:47.40" lane="4" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="359" eventid="19" swimtime="00:01:39.08" lane="2" heatid="19003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="91" birthdate="2012-01-01" gender="M" lastname="Mellenthin" firstname="Linus" license="461669">
              <RESULTS>
                <RESULT resultid="360" eventid="4" swimtime="00:00:49.51" lane="1" heatid="4004" />
                <RESULT resultid="361" eventid="6" swimtime="00:02:11.73" lane="1" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="362" eventid="8" swimtime="00:00:43.43" lane="4" heatid="8003" />
                <RESULT resultid="363" eventid="10" swimtime="00:01:51.10" lane="4" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="364" eventid="18" swimtime="00:00:59.25" lane="2" heatid="18001" />
                <RESULT resultid="365" eventid="20" swimtime="00:01:39.25" lane="1" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="92" birthdate="1997-01-01" gender="M" lastname="Rodriguez Weber" firstname="Adrian" license="171364">
              <RESULTS>
                <RESULT resultid="366" eventid="42" swimtime="00:00:27.16" lane="4" heatid="42008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="93" birthdate="2010-01-01" gender="F" lastname="Schatalin" firstname="Elena" license="435619">
              <RESULTS>
                <RESULT resultid="367" eventid="25" swimtime="00:00:35.25" lane="3" heatid="25009" />
                <RESULT resultid="368" eventid="31" swimtime="00:01:08.47" lane="3" heatid="31009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="369" eventid="33" swimtime="00:01:20.01" lane="3" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="370" eventid="35" swimtime="00:02:50.64" lane="4" heatid="35002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                    <SPLIT distance="150" swimtime="00:02:08.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="371" eventid="41" swimtime="00:00:34.01" lane="2" heatid="41010" />
                <RESULT resultid="372" eventid="43" swimtime="00:00:31.02" lane="3" heatid="43013" />
                <RESULT resultid="373" eventid="47" swimtime="00:01:19.79" lane="1" heatid="47006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="94" birthdate="2009-01-01" gender="M" lastname="Schober" firstname="Florian" license="439713">
              <RESULTS>
                <RESULT resultid="374" eventid="26" swimtime="00:00:34.86" lane="1" heatid="26008" />
                <RESULT resultid="375" eventid="28" swimtime="00:00:35.71" lane="2" heatid="28006" />
                <RESULT resultid="376" eventid="38" swimtime="00:02:58.99" lane="2" heatid="38001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:13.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="377" eventid="42" swimtime="00:00:33.78" lane="1" heatid="42009" />
                <RESULT resultid="378" eventid="44" swimtime="00:00:30.84" lane="4" heatid="44011" />
                <RESULT resultid="379" eventid="46" swimtime="00:01:25.67" lane="3" heatid="46003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="95" birthdate="2003-01-01" gender="M" lastname="Schulze" firstname="Eric" license="298385">
              <RESULTS>
                <RESULT resultid="380" eventid="28" swimtime="00:00:32.31" lane="3" heatid="28009" />
                <RESULT resultid="381" eventid="30" swimtime="00:01:05.42" lane="1" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="382" eventid="34" swimtime="00:01:05.53" lane="4" heatid="34008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="383" eventid="36" swimtime="00:02:36.35" lane="4" heatid="36002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="384" eventid="42" swimtime="00:00:28.42" lane="2" heatid="42007" />
                <RESULT resultid="385" eventid="46" swimtime="00:01:13.28" lane="2" heatid="46006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="386" eventid="54" swimtime="00:02:41.33" lane="4" heatid="54003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:59.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="96" birthdate="2011-01-01" gender="M" lastname="Sommer" firstname="Erik" license="441664">
              <RESULTS>
                <RESULT resultid="387" eventid="4" swimtime="00:00:44.02" lane="3" heatid="4014" />
                <RESULT resultid="388" eventid="8" swimtime="00:00:37.86" lane="4" heatid="8010" />
                <RESULT resultid="389" eventid="10" status="DSQ" swimtime="00:01:40.99" lane="3" heatid="10010" comment="Beim Zielanschlag der Teilstrecke Brust hat der Sportler nicht mit beiden Händen gleichzeitig angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="390" eventid="14" swimtime="00:00:51.96" lane="4" heatid="14010" />
                <RESULT resultid="391" eventid="18" swimtime="00:00:52.75" lane="4" heatid="18012" />
                <RESULT resultid="392" eventid="22" swimtime="00:03:37.59" lane="1" heatid="22002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.83" />
                    <SPLIT distance="100" swimtime="00:01:47.23" />
                    <SPLIT distance="150" swimtime="00:02:52.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="97" birthdate="2005-01-01" gender="M" lastname="Stantke" firstname="Arion" license="344826">
              <RESULTS>
                <RESULT resultid="393" eventid="26" swimtime="00:00:34.34" lane="2" heatid="26004" />
                <RESULT resultid="394" eventid="28" swimtime="00:00:33.87" lane="3" heatid="28005" />
                <RESULT resultid="395" eventid="32" swimtime="00:01:02.26" lane="4" heatid="32006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="396" eventid="42" swimtime="00:00:29.07" lane="3" heatid="42007" />
                <RESULT resultid="397" eventid="44" swimtime="00:00:27.11" lane="2" heatid="44008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="98" birthdate="2007-01-01" gender="M" lastname="Unger" firstname="Tobias" license="404260">
              <RESULTS>
                <RESULT resultid="398" eventid="26" swimtime="00:00:33.02" lane="2" heatid="26003" />
                <RESULT resultid="399" eventid="28" swimtime="00:00:36.68" lane="1" heatid="28003" />
                <RESULT resultid="400" eventid="34" swimtime="00:01:15.31" lane="4" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="401" eventid="42" swimtime="00:00:31.40" lane="1" heatid="42004" />
                <RESULT resultid="402" eventid="44" swimtime="00:00:27.70" lane="4" heatid="44007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="99" birthdate="2009-01-01" gender="F" lastname="Zieb" firstname="Anna Florentine" license="405985">
              <RESULTS>
                <RESULT resultid="403" eventid="29" status="DSQ" swimtime="00:01:20.44" lane="3" heatid="29004" comment="Beim Anschlag an der dritten Wende hat die Sportlerin nicht mit beiden Händen gleichzeitig angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="404" eventid="33" swimtime="00:01:16.05" lane="3" heatid="33008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="405" eventid="41" swimtime="00:00:33.09" lane="3" heatid="41011" />
                <RESULT resultid="406" eventid="43" swimtime="00:00:30.85" lane="4" heatid="43014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100" birthdate="2006-01-01" gender="M" lastname="Zieb" firstname="Tom" license="344952">
              <RESULTS>
                <RESULT resultid="407" eventid="28" swimtime="00:00:35.43" lane="1" heatid="28005" />
                <RESULT resultid="408" eventid="34" swimtime="00:01:12.61" lane="2" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="409" eventid="38" swimtime="00:03:01.31" lane="3" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:27.49" />
                    <SPLIT distance="150" swimtime="00:02:15.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="410" eventid="44" swimtime="00:00:27.86" lane="2" heatid="44007" />
                <RESULT resultid="411" eventid="46" swimtime="00:01:20.76" lane="1" heatid="46005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="412" eventid="54" status="DSQ" swimtime="00:02:46.02" lane="1" heatid="54002" comment="Bei der Wende auf der Teilstrecke Brust hat der Sportler nicht mit beiden Händen gleichzeitig angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:18.82" />
                    <SPLIT distance="150" swimtime="00:02:08.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="309" eventid="11" swimtime="00:02:35.69" lane="1" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                    <SPLIT distance="150" swimtime="00:01:59.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="90" number="1" />
                    <RELAYPOSITION athleteid="96" number="2" />
                    <RELAYPOSITION athleteid="83" number="3" />
                    <RELAYPOSITION athleteid="87" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="310" eventid="23" swimtime="00:02:34.86" lane="4" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:01:25.37" />
                    <SPLIT distance="150" swimtime="00:01:58.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="96" number="1" />
                    <RELAYPOSITION athleteid="86" number="2" />
                    <RELAYPOSITION athleteid="93" number="3" />
                    <RELAYPOSITION athleteid="87" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="311" eventid="40" swimtime="00:01:44.87" lane="4" heatid="40003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.47" />
                    <SPLIT distance="100" swimtime="00:00:52.38" />
                    <SPLIT distance="150" swimtime="00:01:18.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="92" number="1" />
                    <RELAYPOSITION athleteid="100" number="2" />
                    <RELAYPOSITION athleteid="97" number="3" />
                    <RELAYPOSITION athleteid="95" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="312" eventid="40" status="WDR" swimtime="00:00:00.00" lane="1" heatid="40002" />
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="313" eventid="39" swimtime="00:02:06.50" lane="3" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:05.06" />
                    <SPLIT distance="150" swimtime="00:01:36.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="93" number="1" />
                    <RELAYPOSITION athleteid="86" number="2" />
                    <RELAYPOSITION athleteid="84" number="3" />
                    <RELAYPOSITION athleteid="99" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC Freital" nation="GER" region="12" code="3339">
          <ATHLETES>
            <ATHLETE athleteid="214" birthdate="2011-01-01" gender="M" lastname="Börner" firstname="Fynn" license="425572">
              <RESULTS>
                <RESULT resultid="998" eventid="6" swimtime="00:01:36.80" lane="1" heatid="6009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="999" eventid="8" swimtime="00:00:36.21" lane="4" heatid="8019" />
                <RESULT resultid="1000" eventid="14" swimtime="00:00:42.96" lane="1" heatid="14010" />
                <RESULT resultid="1001" eventid="18" swimtime="00:00:44.40" lane="3" heatid="18012" />
                <RESULT resultid="1002" eventid="20" swimtime="00:01:25.86" lane="1" heatid="20015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="215" birthdate="2007-01-01" gender="M" lastname="Feyer" firstname="Luis" license="367868">
              <RESULTS>
                <RESULT resultid="1003" eventid="28" swimtime="00:00:37.18" lane="1" heatid="28002" />
                <RESULT resultid="1004" eventid="32" swimtime="00:01:04.19" lane="3" heatid="32005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1005" eventid="34" swimtime="00:01:15.79" lane="1" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1006" eventid="42" swimtime="00:00:34.03" lane="4" heatid="42003" />
                <RESULT resultid="1007" eventid="44" swimtime="00:00:28.93" lane="2" heatid="44005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="216" birthdate="2010-01-01" gender="F" lastname="Gahner" firstname="Masine" license="406268">
              <RESULTS>
                <RESULT resultid="1008" eventid="25" swimtime="00:00:34.05" lane="2" heatid="25009" />
                <RESULT resultid="1009" eventid="29" swimtime="00:01:19.13" lane="2" heatid="29003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1010" eventid="33" swimtime="00:01:15.28" lane="2" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1011" eventid="43" swimtime="00:00:29.25" lane="2" heatid="43013" />
                <RESULT resultid="1012" eventid="47" swimtime="00:01:15.25" lane="2" heatid="47006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="217" birthdate="2011-01-01" gender="M" lastname="Hentsch" firstname="Oskar René" license="425566">
              <RESULTS>
                <RESULT resultid="1013" eventid="4" swimtime="00:00:42.03" lane="1" heatid="4014" />
                <RESULT resultid="1014" eventid="8" swimtime="00:00:38.88" lane="1" heatid="8007" />
                <RESULT resultid="1015" eventid="10" swimtime="00:01:34.88" lane="1" heatid="10010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1016" eventid="16" swimtime="00:01:31.92" lane="1" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1017" eventid="20" swimtime="00:01:27.07" lane="2" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="218" birthdate="2010-01-01" gender="F" lastname="Heuer" firstname="Lia-Kiara" license="413355">
              <RESULTS>
                <RESULT resultid="1018" eventid="27" swimtime="00:00:42.42" lane="1" heatid="27005" />
                <RESULT resultid="1019" eventid="33" swimtime="00:01:22.97" lane="2" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1020" eventid="41" swimtime="00:00:35.62" lane="1" heatid="41010" />
                <RESULT resultid="1021" eventid="43" swimtime="00:00:31.33" lane="1" heatid="43013" />
                <RESULT resultid="1022" eventid="47" swimtime="00:01:21.76" lane="2" heatid="47002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="219" birthdate="2012-01-01" gender="M" lastname="Kretzschmar" firstname="Nils" license="438792">
              <RESULTS>
                <RESULT resultid="1023" eventid="4" swimtime="00:00:37.20" lane="3" heatid="4013" />
                <RESULT resultid="1024" eventid="8" swimtime="00:00:33.97" lane="3" heatid="8013" />
                <RESULT resultid="1025" eventid="14" swimtime="00:00:40.25" lane="2" heatid="14003" />
                <RESULT resultid="1026" eventid="16" swimtime="00:01:21.57" lane="3" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1027" eventid="20" swimtime="00:01:19.29" lane="3" heatid="20009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="220" birthdate="2009-01-01" gender="F" lastname="Lorenz" firstname="Sophia" license="402585">
              <RESULTS>
                <RESULT resultid="1028" eventid="25" swimtime="00:00:36.21" lane="4" heatid="25006" />
                <RESULT resultid="1029" eventid="33" swimtime="00:01:18.18" lane="3" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1030" eventid="41" swimtime="00:00:35.00" lane="1" heatid="41006" />
                <RESULT resultid="1031" eventid="43" swimtime="00:00:30.92" lane="1" heatid="43010" />
                <RESULT resultid="1032" eventid="47" swimtime="00:01:19.45" lane="4" heatid="47007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="221" birthdate="2010-01-01" gender="F" lastname="Mann" firstname="Emma" license="418262">
              <RESULTS>
                <RESULT resultid="1033" eventid="27" swimtime="00:00:47.41" lane="1" heatid="27001" />
                <RESULT resultid="1034" eventid="31" swimtime="00:01:22.52" lane="4" heatid="31002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1035" eventid="33" status="DSQ" swimtime="00:01:31.18" lane="1" heatid="33001" comment="Die Sportlerin startete vor dem Startsignal">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1036" eventid="43" swimtime="00:00:37.91" lane="2" heatid="43004" />
                <RESULT resultid="1037" eventid="45" swimtime="00:01:45.05" lane="1" heatid="45003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="222" birthdate="2009-01-01" gender="F" lastname="Markert" firstname="Pauline" license="413357">
              <RESULTS>
                <RESULT resultid="1038" eventid="25" swimtime="00:00:38.66" lane="4" heatid="25004" />
                <RESULT resultid="1039" eventid="41" swimtime="00:00:39.72" lane="2" heatid="41003" />
                <RESULT resultid="1040" eventid="43" status="DNS" swimtime="00:00:00.00" lane="2" heatid="43006" />
                <RESULT resultid="1041" eventid="45" swimtime="00:01:33.31" lane="1" heatid="45004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1042" eventid="47" status="DNS" swimtime="00:00:00.00" lane="1" heatid="47004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="223" birthdate="2012-01-01" gender="M" lastname="Matuschka" firstname="Louis" license="452939">
              <RESULTS>
                <RESULT resultid="1043" eventid="6" swimtime="00:01:59.18" lane="2" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1044" eventid="8" swimtime="00:00:47.87" lane="1" heatid="8002" />
                <RESULT resultid="1045" eventid="10" swimtime="00:01:58.50" lane="3" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1046" eventid="18" swimtime="00:00:55.59" lane="2" heatid="18002" />
                <RESULT resultid="1047" eventid="20" swimtime="00:01:49.43" lane="1" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="224" birthdate="2010-01-01" gender="M" lastname="Neubert" firstname="Lino" license="413354">
              <RESULTS>
                <RESULT resultid="1048" eventid="4" swimtime="00:00:40.73" lane="4" heatid="4009" />
                <RESULT resultid="1049" eventid="8" swimtime="00:00:34.02" lane="1" heatid="8013" />
                <RESULT resultid="1050" eventid="10" swimtime="00:01:26.18" lane="2" heatid="10005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1051" eventid="18" swimtime="00:00:44.20" lane="2" heatid="18007" />
                <RESULT resultid="1052" eventid="20" swimtime="00:01:18.03" lane="1" heatid="20010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="225" birthdate="2011-01-01" gender="F" lastname="Neumann" firstname="Antonia" license="429632">
              <RESULTS>
                <RESULT resultid="1053" eventid="3" swimtime="00:00:37.43" lane="1" heatid="3017" />
                <RESULT resultid="1054" eventid="5" swimtime="00:01:29.18" lane="3" heatid="5012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1055" eventid="9" swimtime="00:01:24.77" lane="4" heatid="9010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1056" eventid="17" swimtime="00:00:40.03" lane="3" heatid="17014" />
                <RESULT resultid="1057" eventid="19" swimtime="00:01:14.74" lane="3" heatid="19011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="226" birthdate="2006-01-01" gender="M" lastname="Neumann" firstname="Moritz" license="347128">
              <RESULTS>
                <RESULT resultid="1058" eventid="26" swimtime="00:00:31.66" lane="1" heatid="26005" />
                <RESULT resultid="1059" eventid="36" swimtime="00:02:32.37" lane="1" heatid="36002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="150" swimtime="00:01:54.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1060" eventid="44" swimtime="00:00:27.57" lane="1" heatid="44006" />
                <RESULT resultid="1061" eventid="46" swimtime="00:01:20.61" lane="4" heatid="46005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1062" eventid="48" swimtime="00:01:10.34" lane="1" heatid="48005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="227" birthdate="2007-01-01" gender="M" lastname="Pauer" firstname="Nick" license="367869">
              <RESULTS>
                <RESULT resultid="1063" eventid="28" swimtime="00:00:34.55" lane="1" heatid="28004" />
                <RESULT resultid="1064" eventid="30" swimtime="00:01:19.72" lane="1" heatid="30001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1065" eventid="34" swimtime="00:01:14.09" lane="2" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1066" eventid="42" swimtime="00:00:33.89" lane="1" heatid="42003" />
                <RESULT resultid="1067" eventid="46" swimtime="00:01:19.76" lane="1" heatid="46004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="228" birthdate="2010-01-01" gender="M" lastname="Pink" firstname="Adrian" license="413359">
              <RESULTS>
                <RESULT resultid="1068" eventid="4" swimtime="00:00:36.32" lane="1" heatid="4015" />
                <RESULT resultid="1069" eventid="8" swimtime="00:00:33.37" lane="1" heatid="8014" />
                <RESULT resultid="1070" eventid="10" swimtime="00:01:24.18" lane="3" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1071" eventid="16" swimtime="00:01:20.56" lane="2" heatid="16009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1072" eventid="18" swimtime="00:00:48.04" lane="3" heatid="18006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="229" birthdate="2010-01-01" gender="F" lastname="Röder" firstname="Pauline" license="406267">
              <RESULTS>
                <RESULT resultid="1073" eventid="27" swimtime="00:00:45.97" lane="3" heatid="27001" />
                <RESULT resultid="1074" eventid="33" swimtime="00:01:33.49" lane="1" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1075" eventid="37" swimtime="00:03:38.86" lane="2" heatid="37001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                    <SPLIT distance="100" swimtime="00:01:46.32" />
                    <SPLIT distance="150" swimtime="00:02:44.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1076" eventid="43" swimtime="00:00:38.16" lane="1" heatid="43002" />
                <RESULT resultid="1077" eventid="45" swimtime="00:01:40.50" lane="4" heatid="45003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="230" birthdate="2007-01-01" gender="M" lastname="Rödig" firstname="Luca Maurice" license="362599">
              <RESULTS>
                <RESULT resultid="1078" eventid="26" swimtime="00:00:35.84" lane="4" heatid="26003" />
                <RESULT resultid="1079" eventid="32" swimtime="00:01:06.12" lane="3" heatid="32004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1080" eventid="34" swimtime="00:01:15.10" lane="4" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1081" eventid="42" swimtime="00:00:34.12" lane="2" heatid="42002" />
                <RESULT resultid="1082" eventid="44" swimtime="00:00:28.68" lane="4" heatid="44005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="231" birthdate="1998-01-01" gender="M" lastname="Scharf" firstname="Julien" license="178843">
              <RESULTS>
                <RESULT resultid="1083" eventid="42" swimtime="00:00:32.50" lane="3" heatid="42003" />
                <RESULT resultid="1084" eventid="44" swimtime="00:00:28.73" lane="2" heatid="44006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="232" birthdate="2009-01-01" gender="F" lastname="Schmidt" firstname="Carolyn" license="385998">
              <RESULTS>
                <RESULT resultid="1085" eventid="27" swimtime="00:00:39.38" lane="4" heatid="27006" />
                <RESULT resultid="1086" eventid="31" swimtime="00:01:07.30" lane="3" heatid="31010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1087" eventid="33" swimtime="00:01:17.93" lane="2" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1088" eventid="41" swimtime="00:00:34.22" lane="4" heatid="41011" />
                <RESULT resultid="1089" eventid="43" swimtime="00:00:29.82" lane="1" heatid="43014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="233" birthdate="2006-01-01" gender="M" lastname="Schmidt" firstname="Moritz-Joy" license="347127">
              <RESULTS>
                <RESULT resultid="1090" eventid="28" swimtime="00:00:31.34" lane="1" heatid="28008" />
                <RESULT resultid="1091" eventid="30" status="DSQ" swimtime="00:01:01.37" lane="2" heatid="30003" comment="Beim Anschlag an der dritten Wende hat der Sportler nicht mit beiden Händen gleichzeitig angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1092" eventid="32" swimtime="00:00:55.52" lane="1" heatid="32010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1093" eventid="42" swimtime="00:00:26.80" lane="3" heatid="42011" />
                <RESULT resultid="1094" eventid="44" swimtime="00:00:25.33" lane="1" heatid="44013" />
                <RESULT resultid="2070" eventid="62" swimtime="00:00:31.17" lane="4" heatid="62001" />
                <RESULT resultid="2079" eventid="65" swimtime="00:00:26.83" lane="2" heatid="65001" />
                <RESULT resultid="2098" eventid="69" swimtime="00:00:25.19" lane="1" heatid="69001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="234" birthdate="2011-01-01" gender="M" lastname="Setzer" firstname="Nils" license="425569">
              <RESULTS>
                <RESULT resultid="1095" eventid="6" swimtime="00:01:31.73" lane="3" heatid="6009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1096" eventid="8" swimtime="00:00:33.09" lane="1" heatid="8019" />
                <RESULT resultid="1097" eventid="14" swimtime="00:00:43.53" lane="3" heatid="14010" />
                <RESULT resultid="1098" eventid="18" swimtime="00:00:42.57" lane="2" heatid="18012" />
                <RESULT resultid="1099" eventid="20" swimtime="00:01:16.42" lane="3" heatid="20015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="235" birthdate="2012-01-01" gender="M" lastname="Wiedmann" firstname="Runar" license="448346">
              <RESULTS>
                <RESULT resultid="1100" eventid="4" swimtime="00:00:40.99" lane="1" heatid="4013" />
                <RESULT resultid="1101" eventid="8" swimtime="00:00:34.84" lane="2" heatid="8012" />
                <RESULT resultid="1102" eventid="10" swimtime="00:01:28.02" lane="1" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1103" eventid="16" swimtime="00:01:26.74" lane="3" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1104" eventid="20" swimtime="00:01:19.96" lane="3" heatid="20008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="994" eventid="39" swimtime="00:01:59.27" lane="1" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:00:59.08" />
                    <SPLIT distance="150" swimtime="00:01:28.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="216" number="1" />
                    <RELAYPOSITION athleteid="232" number="2" />
                    <RELAYPOSITION athleteid="220" number="3" />
                    <RELAYPOSITION athleteid="218" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="995" eventid="71" swimtime="00:02:20.12" lane="2" heatid="71002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:50.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="216" number="1" />
                    <RELAYPOSITION athleteid="220" number="2" />
                    <RELAYPOSITION athleteid="218" number="3" />
                    <RELAYPOSITION athleteid="232" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="996" eventid="40" swimtime="00:01:48.55" lane="2" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="100" swimtime="00:00:53.36" />
                    <SPLIT distance="150" swimtime="00:01:20.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="233" number="1" />
                    <RELAYPOSITION athleteid="231" number="2" />
                    <RELAYPOSITION athleteid="226" number="3" />
                    <RELAYPOSITION athleteid="215" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="997" eventid="72" swimtime="00:01:59.13" lane="2" heatid="72002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:04.47" />
                    <SPLIT distance="150" swimtime="00:01:31.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="226" number="1" />
                    <RELAYPOSITION athleteid="227" number="2" />
                    <RELAYPOSITION athleteid="233" number="3" />
                    <RELAYPOSITION athleteid="231" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC Plauen 06" nation="GER" region="12" code="6374">
          <ATHLETES>
            <ATHLETE athleteid="14" birthdate="2006-01-01" gender="F" lastname="Gruber" firstname="Tessa" license="353903">
              <RESULTS>
                <RESULT resultid="52" eventid="25" swimtime="00:00:30.68" lane="3" heatid="25012" />
                <RESULT resultid="53" eventid="27" swimtime="00:00:36.72" lane="2" heatid="27008" />
                <RESULT resultid="54" eventid="35" swimtime="00:02:29.48" lane="3" heatid="35003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="100" swimtime="00:01:14.43" />
                    <SPLIT distance="150" swimtime="00:01:53.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="55" eventid="41" swimtime="00:00:29.40" lane="2" heatid="41013" />
                <RESULT resultid="56" eventid="43" swimtime="00:00:27.67" lane="2" heatid="43016" />
                <RESULT resultid="57" eventid="47" swimtime="00:01:10.31" lane="2" heatid="47009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="58" eventid="53" swimtime="00:02:32.55" lane="2" heatid="53005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:14.58" />
                    <SPLIT distance="150" swimtime="00:01:58.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2044" eventid="56" swimtime="00:00:29.94" lane="4" heatid="56001" />
                <RESULT resultid="2060" eventid="60" swimtime="00:00:34.84" lane="4" heatid="60001" />
                <RESULT resultid="2077" eventid="64" swimtime="00:00:28.58" lane="1" heatid="64001" />
                <RESULT resultid="2093" eventid="68" swimtime="00:00:27.22" lane="1" heatid="68001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="15" birthdate="2012-01-01" gender="F" lastname="Rössel" firstname="Stella" license="439076">
              <RESULTS>
                <RESULT resultid="59" eventid="5" swimtime="00:01:28.65" lane="3" heatid="5011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="60" eventid="9" swimtime="00:01:24.69" lane="1" heatid="9014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="61" eventid="17" swimtime="00:00:39.95" lane="2" heatid="17013" />
                <RESULT resultid="62" eventid="19" swimtime="00:01:15.02" lane="1" heatid="19015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="63" eventid="37" swimtime="00:03:17.91" lane="4" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="150" swimtime="00:02:24.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="64" eventid="51" swimtime="00:02:48.26" lane="4" heatid="51004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:20.72" />
                    <SPLIT distance="150" swimtime="00:02:05.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="ST Erzgebirge" nation="GER" region="12" code="5134">
          <ATHLETES>
            <ATHLETE athleteid="359" birthdate="2012-01-01" gender="M" lastname="Bochmann" firstname="Noa" license="461952">
              <RESULTS>
                <RESULT resultid="1628" eventid="4" swimtime="00:00:50.89" lane="4" heatid="4007" />
                <RESULT resultid="1629" eventid="6" swimtime="00:01:57.00" lane="1" heatid="6004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1630" eventid="8" swimtime="00:00:41.31" lane="3" heatid="8007" />
                <RESULT resultid="1631" eventid="16" status="DSQ" swimtime="00:01:49.07" lane="2" heatid="16001" comment="Der Sportler hat bei der dritten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1632" eventid="18" swimtime="00:00:52.98" lane="2" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="360" birthdate="2011-01-01" gender="M" lastname="Fauska" firstname="Franz" license="458123">
              <RESULTS>
                <RESULT resultid="1633" eventid="4" swimtime="00:00:48.63" lane="4" heatid="4004" />
                <RESULT resultid="1634" eventid="6" swimtime="00:01:48.71" lane="3" heatid="6004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1635" eventid="8" swimtime="00:00:43.95" lane="4" heatid="8006" />
                <RESULT resultid="1636" eventid="18" swimtime="00:00:48.17" lane="1" heatid="18012" />
                <RESULT resultid="1637" eventid="20" swimtime="00:01:42.03" lane="1" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="361" birthdate="2009-01-01" gender="M" lastname="Findeisen" firstname="Erik" license="415866">
              <RESULTS>
                <RESULT resultid="1638" eventid="26" swimtime="00:00:32.89" lane="2" heatid="26008" />
                <RESULT resultid="1639" eventid="28" swimtime="00:00:36.49" lane="3" heatid="28006" />
                <RESULT resultid="1640" eventid="30" swimtime="00:01:11.60" lane="3" heatid="30001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1641" eventid="32" swimtime="00:01:03.28" lane="1" heatid="32008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1642" eventid="34" swimtime="00:01:11.86" lane="2" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1643" eventid="42" swimtime="00:00:30.51" lane="2" heatid="42009" />
                <RESULT resultid="1644" eventid="44" swimtime="00:00:27.80" lane="3" heatid="44011" />
                <RESULT resultid="1645" eventid="46" swimtime="00:01:23.04" lane="1" heatid="46003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1646" eventid="50" swimtime="00:02:52.22" lane="1" heatid="50001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                    <SPLIT distance="150" swimtime="00:02:08.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1647" eventid="54" swimtime="00:02:46.09" lane="2" heatid="54002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:21.20" />
                    <SPLIT distance="150" swimtime="00:02:10.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="362" birthdate="2011-01-01" gender="M" lastname="Frohs" firstname="Erik" license="480943">
              <RESULTS>
                <RESULT resultid="1648" eventid="4" swimtime="00:00:44.86" lane="2" heatid="4006" />
                <RESULT resultid="1649" eventid="6" swimtime="00:02:01.37" lane="3" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1650" eventid="8" swimtime="00:00:37.82" lane="1" heatid="8008" />
                <RESULT resultid="1651" eventid="16" swimtime="00:01:45.92" lane="1" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1652" eventid="18" swimtime="00:00:59.29" lane="3" heatid="18003" />
                <RESULT resultid="1653" eventid="20" swimtime="00:01:36.57" lane="4" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="363" birthdate="2014-01-01" gender="M" lastname="Gläser" firstname="Julian" license="458122">
              <RESULTS>
                <RESULT resultid="1654" eventid="10" swimtime="00:01:51.56" lane="4" heatid="10007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1655" eventid="14" swimtime="00:00:51.45" lane="1" heatid="14007" />
                <RESULT resultid="1656" eventid="18" swimtime="00:01:00.81" lane="1" heatid="18002" />
                <RESULT resultid="1657" eventid="20" swimtime="00:01:48.21" lane="4" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="364" birthdate="2010-01-01" gender="M" lastname="Gläser" firstname="Simon" license="461951">
              <RESULTS>
                <RESULT resultid="1658" eventid="2" swimtime="00:01:40.58" lane="3" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1659" eventid="6" swimtime="00:01:37.52" lane="4" heatid="6010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1660" eventid="8" swimtime="00:00:35.78" lane="1" heatid="8011" />
                <RESULT resultid="1661" eventid="10" swimtime="00:01:32.05" lane="2" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1662" eventid="14" swimtime="00:00:43.04" lane="2" heatid="14005" />
                <RESULT resultid="1663" eventid="18" swimtime="00:00:43.79" lane="3" heatid="18007" />
                <RESULT resultid="1664" eventid="20" swimtime="00:01:24.04" lane="4" heatid="20009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="365" birthdate="2010-01-01" gender="F" lastname="Göhler" firstname="Lucy" license="402479">
              <RESULTS>
                <RESULT resultid="1665" eventid="25" swimtime="00:00:38.37" lane="4" heatid="25009" />
                <RESULT resultid="1666" eventid="29" swimtime="00:01:32.43" lane="3" heatid="29003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1667" eventid="31" swimtime="00:01:15.49" lane="2" heatid="31009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1668" eventid="41" swimtime="00:00:38.60" lane="4" heatid="41010" />
                <RESULT resultid="1669" eventid="43" swimtime="00:00:33.94" lane="4" heatid="43013" />
                <RESULT resultid="1670" eventid="47" swimtime="00:01:25.64" lane="3" heatid="47002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1671" eventid="53" swimtime="00:03:02.40" lane="3" heatid="53001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:28.87" />
                    <SPLIT distance="150" swimtime="00:02:21.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="366" birthdate="2012-01-01" gender="M" lastname="Gottschalk" firstname="Karl" license="461957">
              <RESULTS>
                <RESULT resultid="1672" eventid="4" swimtime="00:00:53.34" lane="2" heatid="4001" />
                <RESULT resultid="1673" eventid="6" swimtime="00:01:54.81" lane="1" heatid="6003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1674" eventid="8" swimtime="00:00:43.52" lane="4" heatid="8004" />
                <RESULT resultid="1675" eventid="18" swimtime="00:00:52.10" lane="1" heatid="18011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="367" birthdate="2008-01-01" gender="M" lastname="Heidenreich" firstname="Luca" license="415867">
              <RESULTS>
                <RESULT resultid="1676" eventid="26" swimtime="00:00:33.37" lane="1" heatid="26004" />
                <RESULT resultid="1677" eventid="28" swimtime="00:00:33.71" lane="2" heatid="28004" />
                <RESULT resultid="1678" eventid="32" swimtime="00:01:07.25" lane="3" heatid="32001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1679" eventid="34" swimtime="00:01:14.03" lane="1" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1680" eventid="38" swimtime="00:02:51.70" lane="1" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                    <SPLIT distance="150" swimtime="00:02:06.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1681" eventid="42" swimtime="00:00:33.18" lane="2" heatid="42003" />
                <RESULT resultid="1682" eventid="44" swimtime="00:00:30.12" lane="3" heatid="44004" />
                <RESULT resultid="1683" eventid="46" swimtime="00:01:20.89" lane="3" heatid="46004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1684" eventid="54" swimtime="00:02:50.91" lane="3" heatid="54002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:22.48" />
                    <SPLIT distance="150" swimtime="00:02:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2065" eventid="61" swimtime="00:00:34.08" lane="4" heatid="61001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="368" birthdate="2007-01-01" gender="F" lastname="Hermann" firstname="Rebekka" license="402476">
              <RESULTS>
                <RESULT resultid="1685" eventid="25" swimtime="00:00:44.71" lane="3" heatid="25002" />
                <RESULT resultid="1686" eventid="31" swimtime="00:01:26.21" lane="1" heatid="31003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1687" eventid="41" swimtime="00:00:41.77" lane="3" heatid="41002" />
                <RESULT resultid="1688" eventid="43" swimtime="00:00:37.63" lane="2" heatid="43002" />
                <RESULT resultid="1689" eventid="47" swimtime="00:01:39.09" lane="1" heatid="47001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="369" birthdate="2011-01-01" gender="F" lastname="Hiemann" firstname="Elisa" license="461993">
              <RESULTS>
                <RESULT resultid="1690" eventid="3" swimtime="00:00:40.39" lane="2" heatid="3008" />
                <RESULT resultid="1691" eventid="5" swimtime="00:01:35.32" lane="2" heatid="5007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1692" eventid="9" swimtime="00:01:27.46" lane="4" heatid="9009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1693" eventid="13" swimtime="00:00:41.18" lane="4" heatid="13010" />
                <RESULT resultid="1694" eventid="15" swimtime="00:01:33.83" lane="4" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1695" eventid="17" swimtime="00:00:42.36" lane="4" heatid="17014" />
                <RESULT resultid="1696" eventid="37" swimtime="00:03:24.87" lane="2" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:41.24" />
                    <SPLIT distance="150" swimtime="00:02:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1697" eventid="51" swimtime="00:03:08.84" lane="2" heatid="51001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:30.55" />
                    <SPLIT distance="150" swimtime="00:02:23.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="370" birthdate="2002-01-01" gender="F" lastname="Katsala" firstname="Mariia" license="458276">
              <RESULTS>
                <RESULT resultid="1698" eventid="25" swimtime="00:00:33.22" lane="4" heatid="25013" />
                <RESULT resultid="1699" eventid="31" swimtime="00:01:04.28" lane="3" heatid="31013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1700" eventid="41" swimtime="00:00:34.18" lane="3" heatid="41007" />
                <RESULT resultid="1701" eventid="43" swimtime="00:00:30.33" lane="1" heatid="43011" />
                <RESULT resultid="1702" eventid="47" swimtime="00:01:12.89" lane="2" heatid="47010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="371" birthdate="2013-01-01" gender="F" lastname="Klaus" firstname="Emma" license="461960">
              <RESULTS>
                <RESULT resultid="1703" eventid="3" swimtime="00:00:49.68" lane="4" heatid="3011" />
                <RESULT resultid="1704" eventid="5" swimtime="00:01:51.39" lane="3" heatid="5004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1705" eventid="7" swimtime="00:00:46.50" lane="4" heatid="7005" />
                <RESULT resultid="1706" eventid="9" swimtime="00:01:53.58" lane="1" heatid="9003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1707" eventid="17" swimtime="00:00:51.01" lane="3" heatid="17007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="372" birthdate="2013-01-01" gender="M" lastname="Konrad" firstname="Christian" license="461953">
              <RESULTS>
                <RESULT resultid="1708" eventid="6" swimtime="00:01:44.47" lane="4" heatid="6005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1709" eventid="8" swimtime="00:00:39.19" lane="4" heatid="8008" />
                <RESULT resultid="1710" eventid="10" swimtime="00:01:41.33" lane="4" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1711" eventid="14" swimtime="00:00:50.93" lane="4" heatid="14004" />
                <RESULT resultid="1712" eventid="18" swimtime="00:00:48.93" lane="3" heatid="18010" />
                <RESULT resultid="1713" eventid="22" swimtime="00:03:43.29" lane="1" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.75" />
                    <SPLIT distance="100" swimtime="00:01:51.98" />
                    <SPLIT distance="150" swimtime="00:02:51.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="373" birthdate="2008-01-01" gender="F" lastname="Künzel" firstname="Collien" license="393376">
              <RESULTS>
                <RESULT resultid="1714" eventid="25" swimtime="00:00:41.01" lane="3" heatid="25003" />
                <RESULT resultid="1715" eventid="31" swimtime="00:01:18.53" lane="1" heatid="31002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1716" eventid="33" swimtime="00:01:31.25" lane="2" heatid="33001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1717" eventid="43" swimtime="00:00:34.07" lane="3" heatid="43004" />
                <RESULT resultid="1718" eventid="47" swimtime="00:01:32.20" lane="1" heatid="47002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="374" birthdate="2012-01-01" gender="F" lastname="Langer" firstname="Mia" license="461959">
              <RESULTS>
                <RESULT resultid="1719" eventid="3" swimtime="00:00:45.93" lane="3" heatid="3006" />
                <RESULT resultid="1720" eventid="7" swimtime="00:00:40.92" lane="4" heatid="7011" />
                <RESULT resultid="1721" eventid="9" swimtime="00:01:48.01" lane="2" heatid="9003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1722" eventid="13" swimtime="00:00:54.01" lane="3" heatid="13003" />
                <RESULT resultid="1723" eventid="17" swimtime="00:00:52.97" lane="1" heatid="17008" />
                <RESULT resultid="1724" eventid="21" swimtime="00:04:00.48" lane="1" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.04" />
                    <SPLIT distance="100" swimtime="00:01:55.94" />
                    <SPLIT distance="150" swimtime="00:03:02.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="375" birthdate="2013-01-01" gender="M" lastname="Langer" firstname="Paul" license="480942">
              <RESULTS>
                <RESULT resultid="1725" eventid="4" swimtime="00:00:57.33" lane="1" heatid="4001" />
                <RESULT resultid="1726" eventid="6" swimtime="00:02:03.42" lane="1" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1727" eventid="8" swimtime="00:00:57.71" lane="1" heatid="8001" />
                <RESULT resultid="1728" eventid="18" swimtime="00:00:55.92" lane="1" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="376" birthdate="2013-01-01" gender="M" lastname="Lehmann" firstname="Jay" license="461955">
              <RESULTS>
                <RESULT resultid="1729" eventid="4" swimtime="00:00:50.43" lane="1" heatid="4002" />
                <RESULT resultid="1730" eventid="8" swimtime="00:00:48.07" lane="2" heatid="8002" />
                <RESULT resultid="1731" eventid="10" swimtime="00:01:54.22" lane="1" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1732" eventid="14" swimtime="00:00:50.73" lane="2" heatid="14002" />
                <RESULT resultid="1733" eventid="20" swimtime="00:01:38.99" lane="3" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1734" eventid="22" swimtime="00:03:59.01" lane="3" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.74" />
                    <SPLIT distance="100" swimtime="00:01:53.77" />
                    <SPLIT distance="150" swimtime="00:03:02.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="377" birthdate="2010-01-01" gender="F" lastname="Lorenz" firstname="Milena" license="417871">
              <RESULTS>
                <RESULT resultid="1735" eventid="25" swimtime="00:00:51.59" lane="3" heatid="25001" />
                <RESULT resultid="1736" eventid="31" swimtime="00:01:35.66" lane="4" heatid="31001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1737" eventid="35" swimtime="00:04:02.17" lane="3" heatid="35001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.40" />
                    <SPLIT distance="100" swimtime="00:01:52.33" />
                    <SPLIT distance="150" swimtime="00:02:57.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1738" eventid="41" swimtime="00:00:45.34" lane="3" heatid="41001" />
                <RESULT resultid="1739" eventid="43" swimtime="00:00:43.22" lane="1" heatid="43001" />
                <RESULT resultid="1740" eventid="51" swimtime="00:03:31.81" lane="1" heatid="51001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:39.39" />
                    <SPLIT distance="150" swimtime="00:02:34.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="378" birthdate="2013-01-01" gender="M" lastname="Meyer" firstname="Sammy" license="458126">
              <RESULTS>
                <RESULT resultid="1741" eventid="4" swimtime="00:00:44.75" lane="1" heatid="4005" />
                <RESULT resultid="1742" eventid="8" swimtime="00:00:37.85" lane="2" heatid="8008" />
                <RESULT resultid="1743" eventid="14" swimtime="00:00:51.32" lane="2" heatid="14001" />
                <RESULT resultid="1744" eventid="16" swimtime="00:01:38.35" lane="1" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1745" eventid="20" swimtime="00:01:30.66" lane="1" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="379" birthdate="2013-01-01" gender="F" lastname="Mildner" firstname="Donna" license="480945">
              <RESULTS>
                <RESULT resultid="1746" eventid="3" swimtime="00:00:56.64" lane="4" heatid="3004" />
                <RESULT resultid="1747" eventid="7" swimtime="00:00:45.92" lane="3" heatid="7001" />
                <RESULT resultid="1748" eventid="13" swimtime="00:01:01.98" lane="1" heatid="13001" />
                <RESULT resultid="1749" eventid="15" swimtime="00:02:04.04" lane="3" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="380" birthdate="2015-01-01" gender="F" lastname="Morgenstern" firstname="Elena" license="471532">
              <RESULTS>
                <RESULT resultid="1750" eventid="3" swimtime="00:00:56.68" lane="2" heatid="3004" />
                <RESULT resultid="1751" eventid="5" swimtime="00:02:00.17" lane="3" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1752" eventid="7" swimtime="00:00:52.02" lane="2" heatid="7003" />
                <RESULT resultid="1753" eventid="15" swimtime="00:02:08.65" lane="4" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1754" eventid="17" swimtime="00:00:54.56" lane="1" heatid="17010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="381" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Annica" license="429663">
              <RESULTS>
                <RESULT resultid="1755" eventid="5" swimtime="00:01:38.13" lane="3" heatid="5007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1756" eventid="7" swimtime="00:00:32.46" lane="4" heatid="7023" />
                <RESULT resultid="1757" eventid="9" swimtime="00:01:25.37" lane="2" heatid="9010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1758" eventid="13" swimtime="00:00:37.53" lane="1" heatid="13010" />
                <RESULT resultid="1759" eventid="17" swimtime="00:00:45.82" lane="3" heatid="17009" />
                <RESULT resultid="1760" eventid="19" swimtime="00:01:14.81" lane="4" heatid="19016">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1761" eventid="37" swimtime="00:03:32.81" lane="3" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                    <SPLIT distance="100" swimtime="00:01:42.60" />
                    <SPLIT distance="150" swimtime="00:02:38.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1762" eventid="51" swimtime="00:02:49.32" lane="3" heatid="51002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:20.29" />
                    <SPLIT distance="150" swimtime="00:02:05.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="382" birthdate="2012-01-01" gender="F" lastname="Müller" firstname="Frieda" license="461992">
              <RESULTS>
                <RESULT resultid="1763" eventid="3" swimtime="00:00:47.10" lane="3" heatid="3013" />
                <RESULT resultid="1764" eventid="5" swimtime="00:01:46.49" lane="3" heatid="5005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1765" eventid="7" swimtime="00:00:36.76" lane="1" heatid="7013" />
                <RESULT resultid="1766" eventid="9" swimtime="00:01:32.89" lane="4" heatid="9008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1767" eventid="15" swimtime="00:01:40.87" lane="1" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1768" eventid="17" swimtime="00:00:50.00" lane="2" heatid="17007" />
                <RESULT resultid="1769" eventid="19" swimtime="00:01:25.45" lane="4" heatid="19009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1770" eventid="37" swimtime="00:03:46.73" lane="3" heatid="37001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.19" />
                    <SPLIT distance="100" swimtime="00:01:47.04" />
                    <SPLIT distance="150" swimtime="00:02:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1771" eventid="51" swimtime="00:03:10.30" lane="3" heatid="51001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:30.27" />
                    <SPLIT distance="150" swimtime="00:02:22.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="383" birthdate="2010-01-01" gender="M" lastname="Neubert" firstname="Alois" license="461950">
              <RESULTS>
                <RESULT resultid="1772" eventid="6" swimtime="00:02:00.09" lane="3" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1773" eventid="8" swimtime="00:00:41.27" lane="4" heatid="8007" />
                <RESULT resultid="1774" eventid="10" swimtime="00:01:50.19" lane="2" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1775" eventid="18" swimtime="00:00:56.55" lane="1" heatid="18003" />
                <RESULT resultid="1776" eventid="20" swimtime="00:01:38.18" lane="4" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="384" birthdate="2009-01-01" gender="M" lastname="Neubert" firstname="Domenic" license="429667">
              <RESULTS>
                <RESULT resultid="1777" eventid="26" swimtime="00:00:36.49" lane="2" heatid="26002" />
                <RESULT resultid="1778" eventid="32" swimtime="00:01:09.92" lane="3" heatid="32002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1779" eventid="34" swimtime="00:01:19.70" lane="4" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1780" eventid="42" status="DSQ" swimtime="00:00:33.69" lane="4" heatid="42009" comment="Der Sportler startete vor dem Startsignal" />
                <RESULT resultid="1781" eventid="44" swimtime="00:00:30.06" lane="2" heatid="44002" />
                <RESULT resultid="1782" eventid="48" swimtime="00:01:24.04" lane="4" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="385" birthdate="2007-01-01" gender="M" lastname="Neubert" firstname="Johannes" license="393375">
              <RESULTS>
                <RESULT resultid="1783" eventid="28" swimtime="00:00:37.18" lane="3" heatid="28002" />
                <RESULT resultid="1784" eventid="32" swimtime="00:01:10.86" lane="4" heatid="32003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1785" eventid="34" swimtime="00:01:20.45" lane="2" heatid="34001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1786" eventid="44" swimtime="00:00:29.66" lane="1" heatid="44004" />
                <RESULT resultid="1787" eventid="46" swimtime="00:01:25.49" lane="3" heatid="46002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1788" eventid="54" swimtime="00:02:48.60" lane="3" heatid="54001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:20.84" />
                    <SPLIT distance="150" swimtime="00:02:10.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="386" birthdate="2011-01-01" gender="F" lastname="Neubert" firstname="Sally" license="429664">
              <RESULTS>
                <RESULT resultid="1789" eventid="3" swimtime="00:00:47.16" lane="1" heatid="3011" />
                <RESULT resultid="1790" eventid="7" swimtime="00:00:42.45" lane="1" heatid="7010" />
                <RESULT resultid="1791" eventid="9" swimtime="00:01:43.14" lane="1" heatid="9005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1792" eventid="13" swimtime="00:00:48.23" lane="2" heatid="13003" />
                <RESULT resultid="1793" eventid="15" swimtime="00:01:43.79" lane="2" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1794" eventid="19" swimtime="00:01:34.33" lane="4" heatid="19007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1795" eventid="35" swimtime="00:03:46.55" lane="1" heatid="35001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.33" />
                    <SPLIT distance="100" swimtime="00:01:46.23" />
                    <SPLIT distance="150" swimtime="00:02:47.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="387" birthdate="2013-01-01" gender="M" lastname="Nordheim" firstname="Matteo" license="461956">
              <RESULTS>
                <RESULT resultid="1796" eventid="4" swimtime="00:01:00.10" lane="3" heatid="4001" />
                <RESULT resultid="1797" eventid="8" swimtime="00:00:47.38" lane="4" heatid="8005" />
                <RESULT resultid="1798" eventid="16" status="DSQ" swimtime="00:02:11.25" lane="3" heatid="16001" comment="Der Sportler hat bei der zweiten und dritten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1799" eventid="20" swimtime="00:01:48.06" lane="2" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="388" birthdate="2013-01-01" gender="F" lastname="Oestreich" firstname="Sophia" license="458275">
              <RESULTS>
                <RESULT resultid="1800" eventid="3" swimtime="00:00:45.89" lane="4" heatid="3012" />
                <RESULT resultid="1801" eventid="7" swimtime="00:00:40.39" lane="3" heatid="7012" />
                <RESULT resultid="1802" eventid="15" swimtime="00:01:44.97" lane="3" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1803" eventid="17" swimtime="00:00:53.69" lane="1" heatid="17004" />
                <RESULT resultid="1804" eventid="19" swimtime="00:01:46.22" lane="4" heatid="19006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="389" birthdate="2015-01-01" gender="F" lastname="Preißler" firstname="Amy" license="480947">
              <RESULTS>
                <RESULT resultid="1805" eventid="3" swimtime="00:01:05.52" lane="3" heatid="3001" />
                <RESULT resultid="1806" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="390" birthdate="1992-01-01" gender="F" lastname="Razeto" firstname="Luisa Marie" license="125894">
              <RESULTS>
                <RESULT resultid="1807" eventid="25" swimtime="00:00:29.99" lane="3" heatid="25013" />
                <RESULT resultid="1808" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="1809" eventid="41" swimtime="00:00:28.41" lane="2" heatid="41014" />
                <RESULT resultid="1810" eventid="43" swimtime="00:00:26.88" lane="2" heatid="43017" />
                <RESULT resultid="2041" eventid="56" swimtime="00:00:29.65" lane="2" heatid="56001" />
                <RESULT resultid="2075" eventid="64" swimtime="00:00:28.30" lane="2" heatid="64001" />
                <RESULT resultid="2091" eventid="68" swimtime="00:00:26.57" lane="2" heatid="68001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="391" birthdate="1986-01-01" gender="M" lastname="Razeto" firstname="Stefano" license="86506">
              <RESULTS>
                <RESULT resultid="1811" eventid="26" swimtime="00:00:26.05" lane="2" heatid="26011" />
                <RESULT resultid="1812" eventid="28" swimtime="00:00:29.51" lane="2" heatid="28009" />
                <RESULT resultid="1813" eventid="42" swimtime="00:00:23.87" lane="2" heatid="42012" />
                <RESULT resultid="1814" eventid="44" swimtime="00:00:22.90" lane="2" heatid="44014" />
                <RESULT resultid="2049" eventid="58" swimtime="00:00:25.44" lane="2" heatid="58001" />
                <RESULT resultid="2067" eventid="62" swimtime="00:00:28.42" lane="2" heatid="62001" />
                <RESULT resultid="2083" eventid="66" swimtime="00:00:23.91" lane="2" heatid="66001" />
                <RESULT resultid="2100" eventid="70" swimtime="00:00:22.24" lane="2" heatid="70001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="392" birthdate="2013-01-01" gender="M" lastname="Rebentrost" firstname="Helios" license="461954">
              <RESULTS>
                <RESULT resultid="1815" eventid="2" swimtime="00:02:12.01" lane="3" heatid="2001">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1816" eventid="4" status="DSQ" swimtime="00:00:48.67" lane="3" heatid="4003" comment="Der Sportler startete vor dem Startsignal" />
                <RESULT resultid="1817" eventid="8" swimtime="00:00:43.44" lane="1" heatid="8003" />
                <RESULT resultid="1818" eventid="14" swimtime="00:00:51.96" lane="4" heatid="14005" />
                <RESULT resultid="1819" eventid="16" swimtime="00:01:48.24" lane="4" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1820" eventid="20" swimtime="00:01:39.60" lane="4" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="393" birthdate="2005-01-01" gender="M" lastname="Reuter" firstname="Erik" license="338774">
              <RESULTS>
                <RESULT resultid="1821" eventid="28" swimtime="00:00:35.99" lane="2" heatid="28003" />
                <RESULT resultid="1822" eventid="32" swimtime="00:00:59.66" lane="4" heatid="32007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1823" eventid="34" swimtime="00:01:10.30" lane="3" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1824" eventid="42" swimtime="00:00:29.93" lane="1" heatid="42006" />
                <RESULT resultid="1825" eventid="44" swimtime="00:00:27.14" lane="3" heatid="44008" />
                <RESULT resultid="1826" eventid="52" swimtime="00:02:18.28" lane="2" heatid="52004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="150" swimtime="00:01:42.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="394" birthdate="2006-01-01" gender="M" lastname="Reuter" firstname="Til" license="382218">
              <RESULTS>
                <RESULT resultid="1827" eventid="28" swimtime="00:00:38.83" lane="4" heatid="28002" />
                <RESULT resultid="1828" eventid="30" swimtime="00:01:19.57" lane="1" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1829" eventid="32" swimtime="00:01:06.66" lane="3" heatid="32003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1830" eventid="42" swimtime="00:00:33.61" lane="3" heatid="42002" />
                <RESULT resultid="1831" eventid="44" swimtime="00:00:29.50" lane="1" heatid="44003" />
                <RESULT resultid="1832" eventid="46" swimtime="00:01:28.66" lane="1" heatid="46002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1833" eventid="50" swimtime="00:03:07.98" lane="4" heatid="50001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:22.78" />
                    <SPLIT distance="150" swimtime="00:02:13.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="395" birthdate="2007-01-01" gender="M" lastname="Richter" firstname="Kimi" license="384061">
              <RESULTS>
                <RESULT resultid="1834" eventid="26" swimtime="00:00:28.72" lane="3" heatid="26009" />
                <RESULT resultid="1835" eventid="28" swimtime="00:00:33.67" lane="1" heatid="28007" />
                <RESULT resultid="1836" eventid="32" swimtime="00:00:57.83" lane="3" heatid="32007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1837" eventid="34" swimtime="00:01:06.09" lane="1" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1838" eventid="44" swimtime="00:00:26.12" lane="1" heatid="44009" />
                <RESULT resultid="1839" eventid="48" swimtime="00:01:07.68" lane="2" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2046" eventid="57" swimtime="00:00:28.99" lane="3" heatid="57001" />
                <RESULT resultid="2064" eventid="61" swimtime="00:00:33.96" lane="1" heatid="61001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="396" birthdate="2002-01-01" gender="F" lastname="Richter" firstname="Nele" license="402475">
              <RESULTS>
                <RESULT resultid="1840" eventid="25" swimtime="00:00:33.05" lane="1" heatid="25013" />
                <RESULT resultid="1841" eventid="29" swimtime="00:01:13.37" lane="3" heatid="29007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1842" eventid="31" swimtime="00:01:05.10" lane="1" heatid="31013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1843" eventid="41" swimtime="00:00:31.20" lane="1" heatid="41014" />
                <RESULT resultid="1844" eventid="43" swimtime="00:00:29.04" lane="1" heatid="43017" />
                <RESULT resultid="1845" eventid="47" swimtime="00:01:13.69" lane="3" heatid="47010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1846" eventid="51" swimtime="00:02:26.36" lane="4" heatid="51005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:07.24" />
                    <SPLIT distance="150" swimtime="00:01:47.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="397" birthdate="2008-01-01" gender="F" lastname="Richter" firstname="Tine" license="429666">
              <RESULTS>
                <RESULT resultid="1847" eventid="25" swimtime="00:00:37.45" lane="1" heatid="25004" />
                <RESULT resultid="1848" eventid="31" swimtime="00:01:10.40" lane="2" heatid="31005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1849" eventid="33" swimtime="00:01:25.00" lane="3" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1850" eventid="41" swimtime="00:00:37.00" lane="3" heatid="41004" />
                <RESULT resultid="1851" eventid="43" swimtime="00:00:31.92" lane="1" heatid="43007" />
                <RESULT resultid="1852" eventid="47" swimtime="00:01:24.32" lane="3" heatid="47003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="398" birthdate="2011-01-01" gender="F" lastname="Rößler" firstname="Lina" license="476556">
              <RESULTS>
                <RESULT resultid="1853" eventid="3" swimtime="00:00:48.35" lane="4" heatid="3010" />
                <RESULT resultid="1854" eventid="7" swimtime="00:00:42.57" lane="4" heatid="7010" />
                <RESULT resultid="1855" eventid="9" swimtime="00:01:51.33" lane="3" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1856" eventid="13" swimtime="00:00:52.41" lane="4" heatid="13003" />
                <RESULT resultid="1857" eventid="17" swimtime="00:00:54.90" lane="3" heatid="17005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="399" birthdate="2007-01-01" gender="F" lastname="Schönherr" firstname="Hannah" license="382221">
              <RESULTS>
                <RESULT resultid="1858" eventid="25" swimtime="00:00:44.15" lane="2" heatid="25002" />
                <RESULT resultid="1859" eventid="29" swimtime="00:01:43.97" lane="4" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1860" eventid="33" swimtime="00:01:38.29" lane="3" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1861" eventid="43" swimtime="00:00:37.57" lane="3" heatid="43002" />
                <RESULT resultid="1862" eventid="47" swimtime="00:01:38.97" lane="3" heatid="47001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1863" eventid="53" swimtime="00:03:36.14" lane="2" heatid="53001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                    <SPLIT distance="100" swimtime="00:01:41.49" />
                    <SPLIT distance="150" swimtime="00:02:46.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="400" birthdate="2011-01-01" gender="F" lastname="Schreiter" firstname="Melissa" license="447078">
              <RESULTS>
                <RESULT resultid="1864" eventid="3" swimtime="00:00:39.17" lane="3" heatid="3016" />
                <RESULT resultid="1865" eventid="5" swimtime="00:01:30.72" lane="1" heatid="5012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1866" eventid="9" swimtime="00:01:23.33" lane="4" heatid="9015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1867" eventid="15" swimtime="00:01:24.71" lane="3" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1868" eventid="17" swimtime="00:00:43.23" lane="2" heatid="17009" />
                <RESULT resultid="1869" eventid="21" swimtime="00:03:01.12" lane="1" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:26.59" />
                    <SPLIT distance="150" swimtime="00:02:16.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1870" eventid="37" swimtime="00:03:12.72" lane="3" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:31.68" />
                    <SPLIT distance="150" swimtime="00:02:22.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1871" eventid="51" swimtime="00:02:53.24" lane="3" heatid="51003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:01:22.77" />
                    <SPLIT distance="150" swimtime="00:02:08.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="401" birthdate="2007-01-01" gender="F" lastname="Steiner" firstname="Tiffany" license="355425">
              <RESULTS>
                <RESULT resultid="1872" eventid="25" swimtime="00:00:35.30" lane="1" heatid="25007" />
                <RESULT resultid="1873" eventid="27" swimtime="00:00:43.37" lane="4" heatid="27004" />
                <RESULT resultid="1874" eventid="33" swimtime="00:01:18.87" lane="1" heatid="33009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1875" eventid="41" swimtime="00:00:35.16" lane="2" heatid="41007" />
                <RESULT resultid="1876" eventid="43" swimtime="00:00:31.87" lane="3" heatid="43008" />
                <RESULT resultid="1877" eventid="51" swimtime="00:02:35.73" lane="3" heatid="51004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:13.87" />
                    <SPLIT distance="150" swimtime="00:01:55.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="402" birthdate="2013-01-01" gender="F" lastname="Stieglitz" firstname="Zoe" license="480944">
              <RESULTS>
                <RESULT resultid="1878" eventid="3" swimtime="00:00:56.32" lane="4" heatid="3002" />
                <RESULT resultid="1879" eventid="7" swimtime="00:00:54.82" lane="3" heatid="7002" />
                <RESULT resultid="1880" eventid="9" status="DSQ" swimtime="00:02:04.07" lane="1" heatid="9001" comment="Beim Zielanschlag der Teilstrecke Brust hat die Sportlerin nicht mit beiden Händen gleichzeitig angeschlagen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1881" eventid="15" swimtime="00:02:14.00" lane="1" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1882" eventid="17" swimtime="00:00:58.66" lane="1" heatid="17001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="403" birthdate="2010-01-01" gender="M" lastname="Treffkorn" firstname="Johann" license="429665">
              <RESULTS>
                <RESULT resultid="1883" eventid="4" status="DNS" swimtime="00:00:00.00" lane="4" heatid="4008" />
                <RESULT resultid="1884" eventid="8" status="DNS" swimtime="00:00:00.00" lane="3" heatid="8006" />
                <RESULT resultid="1885" eventid="14" status="DNS" swimtime="00:00:00.00" lane="3" heatid="14001" />
                <RESULT resultid="1886" eventid="16" status="DNS" swimtime="00:00:00.00" lane="2" heatid="16002" />
                <RESULT resultid="1887" eventid="20" status="DNS" swimtime="00:00:00.00" lane="2" heatid="20003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="404" birthdate="2009-01-01" gender="M" lastname="Tutzschky" firstname="Lukas" license="461949">
              <RESULTS>
                <RESULT resultid="1888" eventid="26" swimtime="00:00:41.53" lane="2" heatid="26001" />
                <RESULT resultid="1889" eventid="32" swimtime="00:01:13.16" lane="2" heatid="32001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1890" eventid="34" status="DSQ" swimtime="00:01:28.59" lane="1" heatid="34001" comment="Der Sportler führte nach der zweiten Wende mit den Beinen wechselseitig Bewegungen aus.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1891" eventid="42" swimtime="00:00:38.85" lane="1" heatid="42001" />
                <RESULT resultid="1892" eventid="44" swimtime="00:00:34.23" lane="3" heatid="44001" />
                <RESULT resultid="1893" eventid="48" swimtime="00:01:35.25" lane="1" heatid="48001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1894" eventid="52" swimtime="00:02:48.01" lane="3" heatid="52001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:23.34" />
                    <SPLIT distance="150" swimtime="00:02:08.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="405" birthdate="2015-01-01" gender="M" lastname="Unger" firstname="Bruno" license="471531">
              <RESULTS>
                <RESULT resultid="1895" eventid="4" swimtime="00:00:51.09" lane="1" heatid="4010" />
                <RESULT resultid="1896" eventid="6" swimtime="00:01:47.83" lane="1" heatid="6006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1897" eventid="8" swimtime="00:00:42.24" lane="1" heatid="8015" />
                <RESULT resultid="1898" eventid="10" swimtime="00:01:46.25" lane="3" heatid="10006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1899" eventid="18" swimtime="00:00:50.68" lane="2" heatid="18008" />
                <RESULT resultid="1900" eventid="20" swimtime="00:01:38.85" lane="1" heatid="20011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="406" birthdate="2014-01-01" gender="F" lastname="Viertel" firstname="Victoria-Luise" license="461991">
              <RESULTS>
                <RESULT resultid="1901" eventid="3" swimtime="00:00:56.90" lane="4" heatid="3007" />
                <RESULT resultid="1902" eventid="5" swimtime="00:02:05.72" lane="1" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1903" eventid="7" swimtime="00:00:54.16" lane="2" heatid="7002" />
                <RESULT resultid="1904" eventid="15" swimtime="00:02:21.31" lane="1" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1905" eventid="17" swimtime="00:00:58.38" lane="2" heatid="17004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="407" birthdate="2006-01-01" gender="F" lastname="Wägner" firstname="Madeleine" license="422523">
              <RESULTS>
                <RESULT resultid="1906" eventid="25" swimtime="00:00:46.24" lane="2" heatid="25001" />
                <RESULT resultid="1907" eventid="27" swimtime="00:00:55.79" lane="4" heatid="27008" />
                <RESULT resultid="1908" eventid="43" swimtime="00:00:40.62" lane="4" heatid="43001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="408" birthdate="2007-01-01" gender="F" lastname="Wanke" firstname="Joy" license="382217">
              <RESULTS>
                <RESULT resultid="1909" eventid="27" status="DNS" swimtime="00:00:00.00" lane="3" heatid="27004" />
                <RESULT resultid="1910" eventid="31" status="DNS" swimtime="00:00:00.00" lane="2" heatid="31001" />
                <RESULT resultid="1911" eventid="33" status="DNS" swimtime="00:00:00.00" lane="4" heatid="33003" />
                <RESULT resultid="1912" eventid="43" status="DNS" swimtime="00:00:00.00" lane="2" heatid="43003" />
                <RESULT resultid="1913" eventid="45" status="DNS" swimtime="00:00:00.00" lane="1" heatid="45002" />
                <RESULT resultid="1914" eventid="53" status="DNS" swimtime="00:00:00.00" lane="1" heatid="53001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="409" birthdate="2005-01-01" gender="M" lastname="Weiß" firstname="Johann" license="327133">
              <RESULTS>
                <RESULT resultid="1915" eventid="26" swimtime="00:00:31.11" lane="1" heatid="26007" />
                <RESULT resultid="1916" eventid="28" swimtime="00:00:33.46" lane="4" heatid="28008" />
                <RESULT resultid="1917" eventid="34" swimtime="00:01:05.99" lane="3" heatid="34007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1918" eventid="42" swimtime="00:00:29.38" lane="4" heatid="42007" />
                <RESULT resultid="1919" eventid="44" swimtime="00:00:27.32" lane="4" heatid="44010" />
                <RESULT resultid="1920" eventid="46" swimtime="00:01:15.42" lane="3" heatid="46005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="410" birthdate="2002-01-01" gender="M" lastname="Weiß" firstname="Konrad" license="298099">
              <RESULTS>
                <RESULT resultid="1921" eventid="28" swimtime="00:00:36.62" lane="4" heatid="28009" />
                <RESULT resultid="1922" eventid="32" swimtime="00:01:07.19" lane="2" heatid="32005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1923" eventid="42" swimtime="00:00:31.20" lane="2" heatid="42005" />
                <RESULT resultid="1924" eventid="44" swimtime="00:00:28.38" lane="3" heatid="44007" />
                <RESULT resultid="1925" eventid="46" status="DNS" swimtime="00:00:00.00" lane="3" heatid="46006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="411" birthdate="2014-01-01" gender="F" lastname="Wilinga" firstname="Joceline" license="480946">
              <RESULTS>
                <RESULT resultid="1926" eventid="3" swimtime="00:01:04.48" lane="2" heatid="3001" />
                <RESULT resultid="1927" eventid="7" status="WDR" swimtime="00:00:00.00" lane="0" heatid="7000" />
                <RESULT resultid="1928" eventid="15" swimtime="00:02:32.48" lane="2" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="412" birthdate="2009-01-01" gender="F" lastname="Wittig" firstname="Emma" license="415865">
              <RESULTS>
                <RESULT resultid="1929" eventid="27" swimtime="00:00:36.21" lane="2" heatid="27006" />
                <RESULT resultid="1930" eventid="29" swimtime="00:01:24.85" lane="1" heatid="29004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1931" eventid="33" swimtime="00:01:18.22" lane="4" heatid="33008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1932" eventid="41" swimtime="00:00:35.13" lane="4" heatid="41007" />
                <RESULT resultid="1933" eventid="43" swimtime="00:00:31.00" lane="2" heatid="43008" />
                <RESULT resultid="1934" eventid="45" swimtime="00:01:21.97" lane="2" heatid="45004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2058" eventid="60" swimtime="00:00:36.42" lane="3" heatid="60001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="417" birthdate="2008-01-01" gender="M" lastname="Kulai" firstname="Vasyl" license="0">
              <RESULTS>
                <RESULT resultid="1950" eventid="26" status="DSQ" swimtime="00:00:36.43" lane="4" heatid="26002" comment="Der Sportler startete vor dem Startsignal" />
                <RESULT resultid="1951" eventid="28" swimtime="00:00:37.63" lane="2" heatid="28005" />
                <RESULT resultid="1952" eventid="32" swimtime="00:01:12.99" lane="4" heatid="32001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1954" eventid="34" swimtime="00:01:22.73" lane="4" heatid="34001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1953" eventid="42" swimtime="00:00:36.75" lane="4" heatid="42001" />
                <RESULT resultid="1955" eventid="44" swimtime="00:00:32.73" lane="4" heatid="44001" />
                <RESULT resultid="1956" eventid="46" swimtime="00:01:25.58" lane="4" heatid="46002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1957" eventid="48" swimtime="00:01:29.48" lane="4" heatid="48001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1614" eventid="40" swimtime="00:01:41.34" lane="3" heatid="40003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.76" />
                    <SPLIT distance="100" swimtime="00:00:52.68" />
                    <SPLIT distance="150" swimtime="00:01:19.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="395" number="1" />
                    <RELAYPOSITION athleteid="393" number="2" />
                    <RELAYPOSITION athleteid="409" number="3" />
                    <RELAYPOSITION athleteid="391" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1615" eventid="72" swimtime="00:01:52.15" lane="3" heatid="72003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                    <SPLIT distance="150" swimtime="00:01:25.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="395" number="1" />
                    <RELAYPOSITION athleteid="409" number="2" />
                    <RELAYPOSITION athleteid="391" number="3" />
                    <RELAYPOSITION athleteid="393" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1616" eventid="39" swimtime="00:01:55.53" lane="2" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                    <SPLIT distance="100" swimtime="00:00:58.67" />
                    <SPLIT distance="150" swimtime="00:01:29.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="370" number="1" />
                    <RELAYPOSITION athleteid="396" number="2" />
                    <RELAYPOSITION athleteid="412" number="3" />
                    <RELAYPOSITION athleteid="390" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1617" eventid="71" swimtime="00:02:07.70" lane="2" heatid="71003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:41.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="370" number="1" />
                    <RELAYPOSITION athleteid="412" number="2" />
                    <RELAYPOSITION athleteid="396" number="3" />
                    <RELAYPOSITION athleteid="390" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1618" eventid="11" swimtime="00:02:18.63" lane="1" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                    <SPLIT distance="150" swimtime="00:01:43.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="381" number="1" />
                    <RELAYPOSITION athleteid="400" number="2" />
                    <RELAYPOSITION athleteid="369" number="3" />
                    <RELAYPOSITION athleteid="364" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1619" eventid="23" swimtime="00:02:33.42" lane="1" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:22.18" />
                    <SPLIT distance="150" swimtime="00:01:59.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="400" number="1" />
                    <RELAYPOSITION athleteid="369" number="2" />
                    <RELAYPOSITION athleteid="381" number="3" />
                    <RELAYPOSITION athleteid="364" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1620" eventid="40" swimtime="00:01:54.65" lane="3" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                    <SPLIT distance="100" swimtime="00:00:55.75" />
                    <SPLIT distance="150" swimtime="00:01:25.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="410" number="1" />
                    <RELAYPOSITION athleteid="361" number="2" />
                    <RELAYPOSITION athleteid="367" number="3" />
                    <RELAYPOSITION athleteid="394" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1621" eventid="72" swimtime="00:02:08.24" lane="3" heatid="72002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:40.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="384" number="1" />
                    <RELAYPOSITION athleteid="367" number="2" />
                    <RELAYPOSITION athleteid="361" number="3" />
                    <RELAYPOSITION athleteid="410" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1622" eventid="39" swimtime="00:02:10.50" lane="1" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                    <SPLIT distance="150" swimtime="00:01:37.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="397" number="1" />
                    <RELAYPOSITION athleteid="381" number="2" />
                    <RELAYPOSITION athleteid="401" number="3" />
                    <RELAYPOSITION athleteid="365" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1623" eventid="71" swimtime="00:02:27.99" lane="3" heatid="71002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:20.46" />
                    <SPLIT distance="150" swimtime="00:01:55.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="397" number="1" />
                    <RELAYPOSITION athleteid="369" number="2" />
                    <RELAYPOSITION athleteid="401" number="3" />
                    <RELAYPOSITION athleteid="381" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1624" eventid="11" swimtime="00:02:34.18" lane="3" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:01:54.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="382" number="1" />
                    <RELAYPOSITION athleteid="362" number="2" />
                    <RELAYPOSITION athleteid="378" number="3" />
                    <RELAYPOSITION athleteid="374" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1625" eventid="23" swimtime="00:02:58.64" lane="2" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                    <SPLIT distance="100" swimtime="00:01:35.37" />
                    <SPLIT distance="150" swimtime="00:02:22.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="362" number="1" />
                    <RELAYPOSITION athleteid="360" number="2" />
                    <RELAYPOSITION athleteid="386" number="3" />
                    <RELAYPOSITION athleteid="382" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1626" eventid="72" swimtime="00:02:22.72" lane="1" heatid="72002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:19.34" />
                    <SPLIT distance="150" swimtime="00:01:53.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="404" number="1" />
                    <RELAYPOSITION athleteid="417" number="2" />
                    <RELAYPOSITION athleteid="394" number="3" />
                    <RELAYPOSITION athleteid="385" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1627" eventid="71" swimtime="00:02:38.54" lane="1" heatid="71002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                    <SPLIT distance="100" swimtime="00:01:22.70" />
                    <SPLIT distance="150" swimtime="00:02:02.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="373" number="1" />
                    <RELAYPOSITION athleteid="400" number="2" />
                    <RELAYPOSITION athleteid="365" number="3" />
                    <RELAYPOSITION athleteid="399" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SV 1919 Grimma" nation="GER" region="12" code="5149">
          <ATHLETES>
            <ATHLETE athleteid="121" birthdate="2015-01-01" gender="F" lastname="Bindheim" firstname="Frieda" license="463477">
              <RESULTS>
                <RESULT resultid="501" eventid="3" swimtime="00:00:54.89" lane="3" heatid="3003" />
                <RESULT resultid="502" eventid="7" swimtime="00:00:53.11" lane="3" heatid="7003" />
                <RESULT resultid="503" eventid="15" swimtime="00:02:00.92" lane="1" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="504" eventid="17" swimtime="00:01:08.32" lane="1" heatid="17002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122" birthdate="2009-01-01" gender="F" lastname="Bindheim" firstname="Lea" license="398054">
              <RESULTS>
                <RESULT resultid="505" eventid="25" swimtime="00:00:38.66" lane="3" heatid="25005" />
                <RESULT resultid="506" eventid="27" swimtime="00:00:49.86" lane="4" heatid="27001" />
                <RESULT resultid="507" eventid="41" swimtime="00:00:41.56" lane="1" heatid="41004" />
                <RESULT resultid="508" eventid="43" swimtime="00:00:35.35" lane="4" heatid="43005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123" birthdate="2009-01-01" gender="M" lastname="Blazy" firstname="Janneck" license="421418">
              <RESULTS>
                <RESULT resultid="509" eventid="26" status="WDR" swimtime="00:00:00.00" lane="0" heatid="26000" />
                <RESULT resultid="510" eventid="28" status="WDR" swimtime="00:00:00.00" lane="0" heatid="28000" />
                <RESULT resultid="511" eventid="32" status="WDR" swimtime="00:00:00.00" lane="0" heatid="32000" />
                <RESULT resultid="512" eventid="34" status="WDR" swimtime="00:00:00.00" lane="0" heatid="34000" />
                <RESULT resultid="513" eventid="42" status="WDR" swimtime="00:00:00.00" lane="0" heatid="42000" />
                <RESULT resultid="514" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
                <RESULT resultid="515" eventid="46" status="WDR" swimtime="00:00:00.00" lane="0" heatid="46000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124" birthdate="2014-01-01" gender="F" lastname="Brauße" firstname="Elena" license="451463">
              <RESULTS>
                <RESULT resultid="516" eventid="3" swimtime="00:00:49.00" lane="2" heatid="3006" />
                <RESULT resultid="517" eventid="5" swimtime="00:01:58.61" lane="2" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="518" eventid="9" swimtime="00:01:51.38" lane="3" heatid="9003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="519" eventid="17" swimtime="00:00:54.54" lane="4" heatid="17005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125" birthdate="2014-01-01" gender="F" lastname="Brendler" firstname="Lena" license="451405">
              <RESULTS>
                <RESULT resultid="520" eventid="3" swimtime="00:00:45.94" lane="1" heatid="3012" />
                <RESULT resultid="521" eventid="7" swimtime="00:00:39.47" lane="3" heatid="7020" />
                <RESULT resultid="522" eventid="9" swimtime="00:01:40.25" lane="1" heatid="9012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="523" eventid="13" swimtime="00:00:48.04" lane="2" heatid="13007" />
                <RESULT resultid="524" eventid="19" swimtime="00:01:33.64" lane="4" heatid="19013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="126" birthdate="2011-01-01" gender="F" lastname="Buchwald" firstname="Mara" license="422685">
              <RESULTS>
                <RESULT resultid="525" eventid="3" swimtime="00:00:35.42" lane="2" heatid="3022" />
                <RESULT resultid="526" eventid="7" swimtime="00:00:33.19" lane="2" heatid="7023" />
                <RESULT resultid="527" eventid="9" swimtime="00:01:27.58" lane="2" heatid="9015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="528" eventid="13" swimtime="00:00:35.37" lane="2" heatid="13010" />
                <RESULT resultid="529" eventid="17" status="DNS" swimtime="00:00:00.00" lane="2" heatid="17014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="127" birthdate="2011-01-01" gender="M" lastname="Dietrich" firstname="Malte" license="422681">
              <RESULTS>
                <RESULT resultid="530" eventid="2" swimtime="00:01:20.24" lane="1" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="531" eventid="4" swimtime="00:00:37.04" lane="2" heatid="4014" />
                <RESULT resultid="532" eventid="8" swimtime="00:00:31.83" lane="2" heatid="8019" />
                <RESULT resultid="533" eventid="14" swimtime="00:00:36.02" lane="2" heatid="14010" />
                <RESULT resultid="534" eventid="16" swimtime="00:01:22.05" lane="2" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="535" eventid="20" swimtime="00:01:12.60" lane="2" heatid="20015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128" birthdate="2015-01-01" gender="F" lastname="Dozsa-Nemeth" firstname="Odett" license="463478">
              <RESULTS>
                <RESULT resultid="536" eventid="3" status="DSQ" swimtime="00:00:46.83" lane="3" heatid="3018" comment="Die Sportlerin hat bei der Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt." />
                <RESULT resultid="537" eventid="5" swimtime="00:02:07.19" lane="2" heatid="5008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="538" eventid="7" swimtime="00:00:43.09" lane="3" heatid="7019" />
                <RESULT resultid="539" eventid="9" swimtime="00:01:54.70" lane="1" heatid="9011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="540" eventid="15" swimtime="00:01:47.04" lane="3" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="541" eventid="19" swimtime="00:01:42.33" lane="3" heatid="19012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129" birthdate="2010-01-01" gender="M" lastname="Duckstein" firstname="Alex" license="412300">
              <RESULTS>
                <RESULT resultid="542" eventid="4" swimtime="00:00:39.04" lane="2" heatid="4009" />
                <RESULT resultid="543" eventid="8" swimtime="00:00:32.32" lane="2" heatid="8013" />
                <RESULT resultid="544" eventid="10" swimtime="00:01:25.15" lane="3" heatid="10005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="545" eventid="16" swimtime="00:01:29.23" lane="4" heatid="16009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="546" eventid="18" swimtime="00:00:45.23" lane="4" heatid="18007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130" birthdate="2011-01-01" gender="F" lastname="Duckstein" firstname="Tanja" license="422686">
              <RESULTS>
                <RESULT resultid="547" eventid="1" swimtime="00:01:22.10" lane="2" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="548" eventid="3" swimtime="00:00:34.33" lane="1" heatid="3022" />
                <RESULT resultid="549" eventid="7" swimtime="00:00:30.73" lane="3" heatid="7023" />
                <RESULT resultid="550" eventid="13" swimtime="00:00:35.12" lane="3" heatid="13010" />
                <RESULT resultid="551" eventid="15" swimtime="00:01:17.40" lane="2" heatid="15014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="552" eventid="19" swimtime="00:01:06.83" lane="2" heatid="19016">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="553" eventid="21" swimtime="00:02:50.75" lane="3" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:18.88" />
                    <SPLIT distance="150" swimtime="00:02:11.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="131" birthdate="2013-01-01" gender="M" lastname="Geleschus" firstname="Yannick" license="449831">
              <RESULTS>
                <RESULT resultid="554" eventid="4" swimtime="00:00:42.53" lane="3" heatid="4007" />
                <RESULT resultid="555" eventid="8" swimtime="00:00:35.97" lane="1" heatid="8009" />
                <RESULT resultid="556" eventid="14" swimtime="00:00:47.93" lane="3" heatid="14004" />
                <RESULT resultid="557" eventid="16" swimtime="00:01:38.24" lane="3" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="558" eventid="20" swimtime="00:01:27.17" lane="3" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="132" birthdate="2015-01-01" gender="F" lastname="Golze" firstname="Clara" license="463479">
              <RESULTS>
                <RESULT resultid="559" eventid="3" status="DNS" swimtime="00:00:00.00" lane="2" heatid="3003" />
                <RESULT resultid="560" eventid="7" status="DNS" swimtime="00:00:00.00" lane="4" heatid="7006" />
                <RESULT resultid="561" eventid="15" status="DNS" swimtime="00:00:00.00" lane="2" heatid="15003" />
                <RESULT resultid="562" eventid="17" status="DNS" swimtime="00:00:00.00" lane="3" heatid="17002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="133" birthdate="2011-01-01" gender="F" lastname="Harbich" firstname="Svea" license="422683">
              <RESULTS>
                <RESULT resultid="563" eventid="5" swimtime="00:01:32.79" lane="4" heatid="5012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="564" eventid="7" swimtime="00:00:33.11" lane="2" heatid="7018" />
                <RESULT resultid="565" eventid="9" swimtime="00:01:25.46" lane="1" heatid="9015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="566" eventid="15" swimtime="00:01:23.16" lane="1" heatid="15014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="567" eventid="17" swimtime="00:00:43.34" lane="1" heatid="17014" />
                <RESULT resultid="568" eventid="19" swimtime="00:01:16.07" lane="1" heatid="19016">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="134" birthdate="2010-01-01" gender="F" lastname="Hartwig" firstname="Annika" license="471349">
              <RESULTS>
                <RESULT resultid="569" eventid="25" swimtime="00:00:44.94" lane="1" heatid="25001" />
                <RESULT resultid="570" eventid="27" swimtime="00:00:44.95" lane="2" heatid="27001" />
                <RESULT resultid="571" eventid="33" swimtime="00:01:32.69" lane="3" heatid="33001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="572" eventid="37" swimtime="00:03:29.83" lane="1" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.51" />
                    <SPLIT distance="100" swimtime="00:01:42.42" />
                    <SPLIT distance="150" swimtime="00:02:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="573" eventid="43" swimtime="00:00:37.32" lane="3" heatid="43001" />
                <RESULT resultid="574" eventid="45" swimtime="00:01:38.09" lane="3" heatid="45003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="135" birthdate="2015-01-01" gender="F" lastname="Hauschild" firstname="Julia" license="463480">
              <RESULTS>
                <RESULT resultid="575" eventid="3" swimtime="00:00:52.81" lane="1" heatid="3003" />
                <RESULT resultid="576" eventid="7" swimtime="00:00:49.91" lane="1" heatid="7004" />
                <RESULT resultid="577" eventid="17" swimtime="00:01:01.07" lane="4" heatid="17003" />
                <RESULT resultid="578" eventid="19" swimtime="00:02:02.57" lane="4" heatid="19012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="136" birthdate="2015-01-01" gender="F" lastname="Heinitz" firstname="Linn" license="467472">
              <RESULTS>
                <RESULT resultid="579" eventid="5" swimtime="00:01:57.87" lane="1" heatid="5008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="580" eventid="7" swimtime="00:00:41.89" lane="1" heatid="7019" />
                <RESULT resultid="581" eventid="9" swimtime="00:01:48.33" lane="3" heatid="9011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="582" eventid="13" swimtime="00:00:50.23" lane="2" heatid="13006" />
                <RESULT resultid="583" eventid="17" swimtime="00:00:53.02" lane="2" heatid="17010" />
                <RESULT resultid="584" eventid="19" swimtime="00:01:39.96" lane="2" heatid="19012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="137" birthdate="2014-01-01" gender="F" lastname="Huerta-Stiehl" firstname="Nelly Johanna" license="451404">
              <RESULTS>
                <RESULT resultid="585" eventid="3" swimtime="00:00:52.21" lane="1" heatid="3007" />
                <RESULT resultid="586" eventid="5" swimtime="00:01:51.87" lane="2" heatid="5009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="587" eventid="15" swimtime="00:01:53.29" lane="3" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="588" eventid="17" swimtime="00:00:50.89" lane="2" heatid="17011" />
                <RESULT resultid="589" eventid="19" swimtime="00:01:41.61" lane="4" heatid="19005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="138" birthdate="2012-01-01" gender="F" lastname="Kobsik" firstname="Zoe" license="449834">
              <RESULTS>
                <RESULT resultid="590" eventid="1" swimtime="00:01:28.61" lane="3" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="591" eventid="7" swimtime="00:00:34.03" lane="1" heatid="7022" />
                <RESULT resultid="592" eventid="9" swimtime="00:01:24.90" lane="3" heatid="9010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="593" eventid="13" swimtime="00:00:37.02" lane="2" heatid="13009" />
                <RESULT resultid="594" eventid="19" swimtime="00:01:14.82" lane="4" heatid="19015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="595" eventid="21" swimtime="00:03:05.76" lane="3" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:29.07" />
                    <SPLIT distance="150" swimtime="00:02:26.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="139" birthdate="2007-01-01" gender="F" lastname="Kösters" firstname="Constanze" license="393103">
              <RESULTS>
                <RESULT resultid="596" eventid="25" swimtime="00:00:35.73" lane="2" heatid="25005" />
                <RESULT resultid="597" eventid="31" swimtime="00:01:10.83" lane="3" heatid="31005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="598" eventid="33" swimtime="00:01:20.56" lane="1" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="599" eventid="41" swimtime="00:00:35.82" lane="3" heatid="41005" />
                <RESULT resultid="600" eventid="47" swimtime="00:01:16.52" lane="3" heatid="47005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="601" eventid="53" swimtime="00:02:54.17" lane="1" heatid="53003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:14.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140" birthdate="2009-01-01" gender="F" lastname="Maneck" firstname="Amilia" license="398061">
              <RESULTS>
                <RESULT resultid="602" eventid="25" swimtime="00:00:32.57" lane="2" heatid="25010" />
                <RESULT resultid="603" eventid="29" swimtime="00:01:16.01" lane="2" heatid="29004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="604" eventid="31" swimtime="00:01:03.52" lane="2" heatid="31010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="605" eventid="41" swimtime="00:00:32.80" lane="2" heatid="41011" />
                <RESULT resultid="606" eventid="43" swimtime="00:00:29.40" lane="3" heatid="43014" />
                <RESULT resultid="607" eventid="47" swimtime="00:01:13.63" lane="2" heatid="47007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="141" birthdate="2007-01-01" gender="M" lastname="Maneck" firstname="Samuel" license="405759">
              <RESULTS>
                <RESULT resultid="608" eventid="26" swimtime="00:00:30.19" lane="3" heatid="26006" />
                <RESULT resultid="609" eventid="28" swimtime="00:00:35.34" lane="4" heatid="28004" />
                <RESULT resultid="610" eventid="30" swimtime="00:01:03.50" lane="3" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="611" eventid="32" swimtime="00:00:57.42" lane="1" heatid="32009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="612" eventid="34" swimtime="00:01:09.13" lane="3" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="613" eventid="42" swimtime="00:00:27.69" lane="3" heatid="42010" />
                <RESULT resultid="614" eventid="44" swimtime="00:00:25.96" lane="4" heatid="44012" />
                <RESULT resultid="615" eventid="48" swimtime="00:01:08.48" lane="4" heatid="48004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2081" eventid="65" swimtime="00:00:27.77" lane="1" heatid="65001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="142" birthdate="2014-01-01" gender="F" lastname="Möbius" firstname="Lotte" license="451461">
              <RESULTS>
                <RESULT resultid="616" eventid="3" status="DSQ" swimtime="00:00:47.99" lane="3" heatid="3009" comment="Die Sportlerin hat bei der Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt." />
                <RESULT resultid="617" eventid="5" swimtime="00:01:55.39" lane="1" heatid="5003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="618" eventid="7" status="DSQ" swimtime="00:00:42.05" lane="1" heatid="7009" comment="Die Sportlerin startete vor dem Startsignal" />
                <RESULT resultid="619" eventid="9" swimtime="00:01:45.71" lane="3" heatid="9004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="620" eventid="17" swimtime="00:00:53.54" lane="4" heatid="17011" />
                <RESULT resultid="621" eventid="19" swimtime="00:01:40.80" lane="2" heatid="19005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143" birthdate="2013-01-01" gender="M" lastname="Munari" firstname="Alessandro" license="445022">
              <RESULTS>
                <RESULT resultid="622" eventid="4" swimtime="00:00:41.01" lane="3" heatid="4012" />
                <RESULT resultid="623" eventid="8" swimtime="00:00:37.11" lane="3" heatid="8011" />
                <RESULT resultid="624" eventid="10" swimtime="00:01:36.61" lane="3" heatid="10004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="625" eventid="16" swimtime="00:01:27.86" lane="1" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="626" eventid="20" swimtime="00:01:21.97" lane="1" heatid="20008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="627" eventid="22" swimtime="00:03:28.79" lane="2" heatid="22002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.38" />
                    <SPLIT distance="100" swimtime="00:01:44.32" />
                    <SPLIT distance="150" swimtime="00:02:47.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144" birthdate="2015-01-01" gender="F" lastname="Naumann" firstname="Phyllis Maira" license="463481">
              <RESULTS>
                <RESULT resultid="628" eventid="3" swimtime="00:00:59.76" lane="4" heatid="3003" />
                <RESULT resultid="629" eventid="7" swimtime="00:00:50.34" lane="2" heatid="7004" />
                <RESULT resultid="630" eventid="17" swimtime="00:01:02.04" lane="2" heatid="17002" />
                <RESULT resultid="631" eventid="19" swimtime="00:01:51.94" lane="2" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145" birthdate="2006-01-01" gender="M" lastname="Oelschläger" firstname="Jake" license="355390">
              <RESULTS>
                <RESULT resultid="632" eventid="26" swimtime="00:00:28.97" lane="3" heatid="26010" />
                <RESULT resultid="633" eventid="30" swimtime="00:01:05.47" lane="3" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="634" eventid="32" swimtime="00:00:56.72" lane="3" heatid="32010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="635" eventid="34" swimtime="00:01:07.20" lane="1" heatid="34007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="636" eventid="42" swimtime="00:00:27.31" lane="2" heatid="42011" />
                <RESULT resultid="637" eventid="44" swimtime="00:00:24.82" lane="2" heatid="44013" />
                <RESULT resultid="638" eventid="48" swimtime="00:01:06.86" lane="3" heatid="48005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2047" eventid="57" swimtime="00:00:28.79" lane="1" heatid="57001" />
                <RESULT resultid="2080" eventid="65" swimtime="00:00:27.22" lane="3" heatid="65001" />
                <RESULT resultid="2097" eventid="69" swimtime="00:00:24.98" lane="3" heatid="69001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="146" birthdate="2015-01-01" gender="F" lastname="Otto" firstname="Pia" license="463476">
              <RESULTS>
                <RESULT resultid="639" eventid="3" swimtime="00:00:46.04" lane="2" heatid="3018" />
                <RESULT resultid="640" eventid="5" swimtime="00:01:57.38" lane="3" heatid="5008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="641" eventid="7" swimtime="00:00:44.15" lane="2" heatid="7019" />
                <RESULT resultid="642" eventid="9" swimtime="00:01:48.32" lane="2" heatid="9011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="643" eventid="13" swimtime="00:00:56.08" lane="3" heatid="13006" />
                <RESULT resultid="644" eventid="15" status="DSQ" swimtime="00:01:42.87" lane="2" heatid="15010" comment="Die Sportlerin hat bei der dritten Wende nach Verlassen der Rückenlage nicht unverzüglich die eigentliche Wendenbewegung ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147" birthdate="2015-01-01" gender="F" lastname="Päßler" firstname="Emma" license="463482">
              <RESULTS>
                <RESULT resultid="645" eventid="3" swimtime="00:00:57.52" lane="2" heatid="3002" />
                <RESULT resultid="646" eventid="7" swimtime="00:00:47.95" lane="3" heatid="7004" />
                <RESULT resultid="647" eventid="15" swimtime="00:02:07.25" lane="2" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="648" eventid="19" swimtime="00:01:55.33" lane="1" heatid="19012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="148" birthdate="2014-01-01" gender="M" lastname="Polzin" firstname="Franz" license="451411">
              <RESULTS>
                <RESULT resultid="649" eventid="4" swimtime="00:00:45.60" lane="1" heatid="4006" />
                <RESULT resultid="650" eventid="8" swimtime="00:00:42.03" lane="2" heatid="8007" />
                <RESULT resultid="651" eventid="10" swimtime="00:01:42.11" lane="2" heatid="10007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="652" eventid="16" swimtime="00:01:41.18" lane="4" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="653" eventid="18" swimtime="00:00:56.99" lane="4" heatid="18003" />
                <RESULT resultid="654" eventid="20" swimtime="00:01:35.37" lane="1" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149" birthdate="2004-01-01" gender="M" lastname="Polzin" firstname="Paul" license="277805">
              <RESULTS>
                <RESULT resultid="655" eventid="26" swimtime="00:00:28.71" lane="2" heatid="26007" />
                <RESULT resultid="656" eventid="30" swimtime="00:01:05.43" lane="3" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="657" eventid="32" swimtime="00:00:59.18" lane="3" heatid="32011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="658" eventid="34" swimtime="00:01:07.39" lane="1" heatid="34008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="659" eventid="42" swimtime="00:00:28.16" lane="4" heatid="42012" />
                <RESULT resultid="660" eventid="44" swimtime="00:00:27.76" lane="4" heatid="44014" />
                <RESULT resultid="661" eventid="48" swimtime="00:01:08.22" lane="1" heatid="48006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150" birthdate="2009-01-01" gender="F" lastname="Rasmussen" firstname="Helen" license="398058">
              <RESULTS>
                <RESULT resultid="662" eventid="31" swimtime="00:01:11.33" lane="4" heatid="31010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="663" eventid="33" swimtime="00:01:24.10" lane="2" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="664" eventid="41" swimtime="00:00:36.54" lane="1" heatid="41007" />
                <RESULT resultid="665" eventid="43" swimtime="00:00:31.58" lane="3" heatid="43009" />
                <RESULT resultid="666" eventid="47" swimtime="00:01:25.92" lane="4" heatid="47004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="151" birthdate="2008-01-01" gender="F" lastname="Säbisch" firstname="Kyra" license="389131">
              <RESULTS>
                <RESULT resultid="667" eventid="25" swimtime="00:00:33.09" lane="1" heatid="25011" />
                <RESULT resultid="668" eventid="27" swimtime="00:00:37.53" lane="2" heatid="27007" />
                <RESULT resultid="669" eventid="41" swimtime="00:00:31.81" lane="3" heatid="41012" />
                <RESULT resultid="670" eventid="43" swimtime="00:00:29.80" lane="2" heatid="43012" />
                <RESULT resultid="2054" eventid="59" swimtime="00:00:36.73" lane="3" heatid="59001" />
                <RESULT resultid="2074" eventid="63" swimtime="00:00:31.43" lane="4" heatid="63001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="152" birthdate="2015-01-01" gender="M" lastname="Schewelew" firstname="Egor" license="463483">
              <RESULTS>
                <RESULT resultid="671" eventid="4" swimtime="00:00:49.26" lane="3" heatid="4010" />
                <RESULT resultid="672" eventid="8" swimtime="00:00:44.50" lane="3" heatid="8015" />
                <RESULT resultid="673" eventid="10" swimtime="00:01:55.17" lane="2" heatid="10006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="674" eventid="16" swimtime="00:01:51.71" lane="1" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="675" eventid="18" swimtime="00:01:01.34" lane="3" heatid="18008" />
                <RESULT resultid="676" eventid="20" swimtime="00:01:43.73" lane="3" heatid="20011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="153" birthdate="2008-01-01" gender="M" lastname="Schmutzer" firstname="Domenik" license="398057">
              <RESULTS>
                <RESULT resultid="677" eventid="26" swimtime="00:00:31.17" lane="4" heatid="26006" />
                <RESULT resultid="678" eventid="28" swimtime="00:00:32.91" lane="2" heatid="28007" />
                <RESULT resultid="679" eventid="32" swimtime="00:00:59.18" lane="1" heatid="32007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="680" eventid="38" swimtime="00:02:44.56" lane="3" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:15.61" />
                    <SPLIT distance="150" swimtime="00:02:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="681" eventid="42" swimtime="00:00:31.63" lane="4" heatid="42005" />
                <RESULT resultid="682" eventid="44" swimtime="00:00:26.43" lane="1" heatid="44010" />
                <RESULT resultid="683" eventid="46" swimtime="00:01:13.55" lane="2" heatid="46004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="684" eventid="54" swimtime="00:02:35.31" lane="1" heatid="54003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                    <SPLIT distance="100" swimtime="00:01:13.73" />
                    <SPLIT distance="150" swimtime="00:01:58.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2062" eventid="61" swimtime="00:00:32.92" lane="2" heatid="61001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154" birthdate="2014-01-01" gender="F" lastname="Seemann" firstname="Emma" license="451406">
              <RESULTS>
                <RESULT resultid="685" eventid="3" swimtime="00:00:48.85" lane="3" heatid="3011" />
                <RESULT resultid="686" eventid="5" swimtime="00:01:57.64" lane="4" heatid="5009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="687" eventid="7" swimtime="00:00:41.02" lane="4" heatid="7020" />
                <RESULT resultid="688" eventid="15" swimtime="00:01:50.37" lane="2" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="689" eventid="17" swimtime="00:00:50.68" lane="1" heatid="17011" />
                <RESULT resultid="690" eventid="19" swimtime="00:01:35.63" lane="1" heatid="19007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="155" birthdate="2013-01-01" gender="F" lastname="Sehr" firstname="Liska Amelia" license="444105">
              <RESULTS>
                <RESULT resultid="691" eventid="3" swimtime="00:00:46.64" lane="2" heatid="3010" />
                <RESULT resultid="692" eventid="5" swimtime="00:01:48.88" lane="4" heatid="5010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="693" eventid="9" status="DSQ" swimtime="00:01:40.42" lane="2" heatid="9006" comment="Die Sportlerin startete vor dem Startsignal">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="694" eventid="17" swimtime="00:00:49.80" lane="1" heatid="17012" />
                <RESULT resultid="695" eventid="19" swimtime="00:01:32.91" lane="3" heatid="19006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156" birthdate="2012-01-01" gender="M" lastname="Stäudte" firstname="Vincent" license="436853">
              <RESULTS>
                <RESULT resultid="696" eventid="2" swimtime="00:01:21.51" lane="1" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="697" eventid="4" swimtime="00:00:34.41" lane="2" heatid="4013" />
                <RESULT resultid="698" eventid="8" swimtime="00:00:31.81" lane="2" heatid="8018" />
                <RESULT resultid="699" eventid="10" swimtime="00:01:17.65" lane="2" heatid="10009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="700" eventid="14" swimtime="00:00:36.04" lane="3" heatid="14009" />
                <RESULT resultid="701" eventid="16" swimtime="00:01:15.42" lane="2" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="702" eventid="20" swimtime="00:01:11.24" lane="3" heatid="20014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="703" eventid="22" swimtime="00:02:51.23" lane="3" heatid="22003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:19.57" />
                    <SPLIT distance="150" swimtime="00:02:10.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157" birthdate="2014-01-01" gender="F" lastname="Streubel" firstname="Eliana Malea" license="451402">
              <RESULTS>
                <RESULT resultid="704" eventid="3" swimtime="00:00:49.93" lane="3" heatid="3007" />
                <RESULT resultid="705" eventid="5" swimtime="00:01:58.49" lane="1" heatid="5009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="706" eventid="7" swimtime="00:00:42.72" lane="2" heatid="7006" />
                <RESULT resultid="707" eventid="15" status="DSQ" swimtime="00:01:51.57" lane="1" heatid="15004" comment="Die Sportlerin hat auf der dritten Teilstrecke die Schwimmlage verlassen.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="708" eventid="17" swimtime="00:00:53.30" lane="3" heatid="17004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="158" birthdate="2013-01-01" gender="M" lastname="Thiele" firstname="Henrik" license="451456">
              <RESULTS>
                <RESULT resultid="709" eventid="4" swimtime="00:00:43.20" lane="2" heatid="4007" />
                <RESULT resultid="710" eventid="6" swimtime="00:01:46.72" lane="4" heatid="6007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="711" eventid="8" swimtime="00:00:36.65" lane="4" heatid="8017" />
                <RESULT resultid="712" eventid="10" swimtime="00:01:36.71" lane="4" heatid="10004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="713" eventid="14" swimtime="00:00:46.36" lane="1" heatid="14004" />
                <RESULT resultid="714" eventid="18" swimtime="00:00:47.32" lane="1" heatid="18006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="159" birthdate="2013-01-01" gender="F" lastname="Voigt" firstname="Sophia" license="444104">
              <RESULTS>
                <RESULT resultid="715" eventid="3" swimtime="00:00:38.86" lane="3" heatid="3020" />
                <RESULT resultid="716" eventid="7" swimtime="00:00:33.72" lane="2" heatid="7021" />
                <RESULT resultid="717" eventid="13" swimtime="00:00:44.66" lane="3" heatid="13008" />
                <RESULT resultid="718" eventid="15" swimtime="00:01:25.77" lane="2" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="719" eventid="19" swimtime="00:01:16.83" lane="2" heatid="19014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="720" eventid="21" swimtime="00:03:25.17" lane="3" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                    <SPLIT distance="100" swimtime="00:01:38.68" />
                    <SPLIT distance="150" swimtime="00:02:41.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2012-01-01" gender="F" lastname="Wandschneider" firstname="Marie" license="436844">
              <RESULTS>
                <RESULT resultid="721" eventid="3" swimtime="00:00:42.33" lane="3" heatid="3014" />
                <RESULT resultid="722" eventid="7" swimtime="00:00:38.62" lane="1" heatid="7014" />
                <RESULT resultid="723" eventid="13" swimtime="00:00:45.20" lane="4" heatid="13004" />
                <RESULT resultid="724" eventid="15" swimtime="00:01:33.47" lane="4" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="725" eventid="19" swimtime="00:01:29.01" lane="3" heatid="19008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2011-01-01" gender="F" lastname="Wilhelm" firstname="Linda" license="436850">
              <RESULTS>
                <RESULT resultid="726" eventid="3" swimtime="00:00:42.07" lane="3" heatid="3017" />
                <RESULT resultid="727" eventid="5" swimtime="00:01:42.73" lane="1" heatid="5006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="728" eventid="7" swimtime="00:00:35.62" lane="3" heatid="7016" />
                <RESULT resultid="729" eventid="15" swimtime="00:01:29.91" lane="4" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="730" eventid="17" swimtime="00:00:48.04" lane="2" heatid="17008" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="495" eventid="11" swimtime="00:02:04.66" lane="2" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:01.84" />
                    <SPLIT distance="150" swimtime="00:01:32.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="156" number="1" />
                    <RELAYPOSITION athleteid="130" number="2" />
                    <RELAYPOSITION athleteid="127" number="3" />
                    <RELAYPOSITION athleteid="129" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="496" eventid="23" swimtime="00:02:22.10" lane="2" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                    <SPLIT distance="150" swimtime="00:01:51.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="156" number="1" />
                    <RELAYPOSITION athleteid="133" number="2" />
                    <RELAYPOSITION athleteid="126" number="3" />
                    <RELAYPOSITION athleteid="130" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="497" eventid="39" swimtime="00:01:59.51" lane="3" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                    <SPLIT distance="100" swimtime="00:00:58.69" />
                    <SPLIT distance="150" swimtime="00:01:29.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="140" number="1" />
                    <RELAYPOSITION athleteid="130" number="2" />
                    <RELAYPOSITION athleteid="150" number="3" />
                    <RELAYPOSITION athleteid="151" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="499" eventid="71" swimtime="00:02:14.86" lane="3" heatid="71003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:44.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="139" number="1" />
                    <RELAYPOSITION athleteid="151" number="2" />
                    <RELAYPOSITION athleteid="140" number="3" />
                    <RELAYPOSITION athleteid="150" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="498" eventid="40" swimtime="00:01:41.62" lane="2" heatid="40003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.98" />
                    <SPLIT distance="100" swimtime="00:00:50.07" />
                    <SPLIT distance="150" swimtime="00:01:15.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="145" number="1" />
                    <RELAYPOSITION athleteid="141" number="2" />
                    <RELAYPOSITION athleteid="149" number="3" />
                    <RELAYPOSITION athleteid="153" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="500" eventid="72" swimtime="00:01:53.94" lane="2" heatid="72003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="100" swimtime="00:01:01.47" />
                    <SPLIT distance="150" swimtime="00:01:29.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="149" number="1" />
                    <RELAYPOSITION athleteid="153" number="2" />
                    <RELAYPOSITION athleteid="141" number="3" />
                    <RELAYPOSITION athleteid="145" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SV 1990 Zschopau" nation="GER" region="12" code="3382">
          <ATHLETES>
            <ATHLETE athleteid="162" birthdate="2013-01-01" gender="F" lastname="Decker" firstname="Helene" license="464574">
              <RESULTS>
                <RESULT resultid="731" eventid="3" swimtime="00:00:50.62" lane="1" heatid="3008" />
                <RESULT resultid="732" eventid="5" swimtime="00:01:58.98" lane="1" heatid="5004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="733" eventid="9" swimtime="00:01:48.38" lane="3" heatid="9006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="734" eventid="17" swimtime="00:00:56.10" lane="1" heatid="17006" />
                <RESULT resultid="735" eventid="19" swimtime="00:01:34.00" lane="1" heatid="19006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163" birthdate="2009-01-01" gender="M" lastname="Hildermann" firstname="Conner" license="477581">
              <RESULTS>
                <RESULT resultid="736" eventid="26" swimtime="00:00:41.38" lane="3" heatid="26001" />
                <RESULT resultid="737" eventid="28" swimtime="00:00:47.44" lane="1" heatid="28001" />
                <RESULT resultid="738" eventid="32" swimtime="00:01:31.92" lane="1" heatid="32001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="739" eventid="44" swimtime="00:00:39.31" lane="1" heatid="44001" />
                <RESULT resultid="740" eventid="46" swimtime="00:01:46.49" lane="3" heatid="46001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164" birthdate="2009-01-01" gender="F" lastname="Hunger" firstname="Lea" license="402166">
              <RESULTS>
                <RESULT resultid="741" eventid="25" swimtime="00:00:34.16" lane="1" heatid="25010" />
                <RESULT resultid="742" eventid="27" swimtime="00:00:39.08" lane="1" heatid="27006" />
                <RESULT resultid="743" eventid="33" swimtime="00:01:18.33" lane="1" heatid="33008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="744" eventid="41" swimtime="00:00:34.03" lane="2" heatid="41006" />
                <RESULT resultid="745" eventid="45" swimtime="00:01:29.45" lane="3" heatid="45004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="746" eventid="47" swimtime="00:01:17.88" lane="1" heatid="47007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165" birthdate="2013-01-01" gender="F" lastname="Keller" firstname="Emma" license="460563">
              <RESULTS>
                <RESULT resultid="747" eventid="3" swimtime="00:00:45.00" lane="1" heatid="3013" />
                <RESULT resultid="748" eventid="7" swimtime="00:00:37.85" lane="2" heatid="7013" />
                <RESULT resultid="749" eventid="13" swimtime="00:00:45.48" lane="1" heatid="13008" />
                <RESULT resultid="750" eventid="19" swimtime="00:01:26.88" lane="1" heatid="19014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="751" eventid="21" swimtime="00:03:33.56" lane="3" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                    <SPLIT distance="100" swimtime="00:01:41.47" />
                    <SPLIT distance="150" swimtime="00:02:44.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166" birthdate="2006-01-01" gender="F" lastname="Kreißig" firstname="Lilly" license="393190">
              <RESULTS>
                <RESULT resultid="752" eventid="25" swimtime="00:00:35.61" lane="1" heatid="25012" />
                <RESULT resultid="753" eventid="29" swimtime="00:01:15.64" lane="1" heatid="29006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="754" eventid="33" swimtime="00:01:17.22" lane="1" heatid="33010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="755" eventid="41" swimtime="00:00:33.22" lane="1" heatid="41013" />
                <RESULT resultid="756" eventid="49" swimtime="00:02:59.27" lane="2" heatid="49001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:21.52" />
                    <SPLIT distance="150" swimtime="00:02:10.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="757" eventid="53" swimtime="00:02:51.30" lane="1" heatid="53004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:21.05" />
                    <SPLIT distance="150" swimtime="00:02:11.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="2014-01-01" gender="F" lastname="Meusel" firstname="Lotta Chayenne" license="474377">
              <RESULTS>
                <RESULT resultid="758" eventid="3" swimtime="00:00:54.39" lane="2" heatid="3005" />
                <RESULT resultid="759" eventid="7" swimtime="00:00:49.44" lane="2" heatid="7005" />
                <RESULT resultid="760" eventid="17" swimtime="00:00:58.91" lane="4" heatid="17004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="168" birthdate="2008-01-01" gender="M" lastname="Meusel" firstname="Noah Joel" license="393191">
              <RESULTS>
                <RESULT resultid="761" eventid="32" swimtime="00:01:04.67" lane="4" heatid="32005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="762" eventid="42" swimtime="00:00:31.91" lane="4" heatid="42004" />
                <RESULT resultid="763" eventid="44" swimtime="00:00:28.75" lane="1" heatid="44005" />
                <RESULT resultid="764" eventid="52" swimtime="00:02:27.65" lane="2" heatid="52003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:50.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169" birthdate="2014-01-01" gender="M" lastname="Reuter" firstname="Nils" license="464573">
              <RESULTS>
                <RESULT resultid="765" eventid="4" status="DSQ" swimtime="00:00:47.73" lane="4" heatid="4005" comment="Bei der Wende hat der Sportler die Wand verlassen, bevor die Rückenlage eingenommen war." />
                <RESULT resultid="766" eventid="8" swimtime="00:00:41.12" lane="2" heatid="8006" />
                <RESULT resultid="767" eventid="10" swimtime="00:01:43.26" lane="1" heatid="10007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="768" eventid="14" swimtime="00:00:52.65" lane="1" heatid="14003" />
                <RESULT resultid="769" eventid="18" swimtime="00:00:57.24" lane="3" heatid="18009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170" birthdate="2012-01-01" gender="F" lastname="Ruprecht" firstname="Sarina Svenja" license="478743">
              <RESULTS>
                <RESULT resultid="770" eventid="3" swimtime="00:00:56.28" lane="1" heatid="3005" />
                <RESULT resultid="771" eventid="5" swimtime="00:01:53.21" lane="3" heatid="5003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="772" eventid="17" swimtime="00:00:53.66" lane="4" heatid="17006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="171" birthdate="2010-01-01" gender="M" lastname="Zingler" firstname="Gustav Albert" license="409207">
              <RESULTS>
                <RESULT resultid="773" eventid="6" swimtime="00:01:17.65" lane="2" heatid="6010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="774" eventid="8" swimtime="00:00:27.59" lane="2" heatid="8020" />
                <RESULT resultid="775" eventid="10" swimtime="00:01:12.37" lane="2" heatid="10011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="776" eventid="14" swimtime="00:00:30.02" lane="2" heatid="14011" />
                <RESULT resultid="777" eventid="18" swimtime="00:00:34.61" lane="2" heatid="18013" />
                <RESULT resultid="778" eventid="20" swimtime="00:01:03.28" lane="2" heatid="20016">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172" birthdate="2007-01-01" gender="F" lastname="Zingler" firstname="Lotte Pauline" license="365814">
              <RESULTS>
                <RESULT resultid="779" eventid="25" swimtime="00:00:34.96" lane="2" heatid="25007" />
                <RESULT resultid="780" eventid="29" swimtime="00:01:20.01" lane="1" heatid="29002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="781" eventid="43" swimtime="00:00:31.77" lane="2" heatid="43009" />
                <RESULT resultid="782" eventid="47" swimtime="00:01:16.37" lane="2" heatid="47005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1958" eventid="11" swimtime="00:02:26.72" lane="4" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:18.32" />
                    <SPLIT distance="150" swimtime="00:01:59.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="165" number="1" />
                    <RELAYPOSITION athleteid="162" number="2" />
                    <RELAYPOSITION athleteid="169" number="3" />
                    <RELAYPOSITION athleteid="171" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SV Fortschritt Pirna" nation="GER" region="12" code="3387">
          <ATHLETES>
            <ATHLETE athleteid="4" birthdate="2012-01-01" gender="M" lastname="Adler" firstname="Bendix" license="448850">
              <RESULTS>
                <RESULT resultid="20" eventid="6" swimtime="00:01:24.39" lane="2" heatid="6008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="21" eventid="10" swimtime="00:01:18.79" lane="1" heatid="10009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="22" eventid="18" swimtime="00:00:38.66" lane="2" heatid="18011" />
                <RESULT resultid="23" eventid="22" status="DSQ" swimtime="00:02:53.53" lane="1" heatid="22003" comment="Der Sportler führte während der Teilstrecke Schmetterling, nach dem Start und bei der Wende mehrere Brustbeinschläge aus.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                    <SPLIT distance="150" swimtime="00:02:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="24" eventid="38" swimtime="00:03:01.93" lane="4" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:28.46" />
                    <SPLIT distance="150" swimtime="00:02:16.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="25" eventid="52" swimtime="00:02:37.42" lane="3" heatid="52002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:01:16.12" />
                    <SPLIT distance="150" swimtime="00:01:58.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Schneeberg Schwimmen" nation="GER" region="12" code="7124">
          <ATHLETES>
            <ATHLETE athleteid="343" birthdate="2011-01-01" gender="M" lastname="Güßmann" firstname="Ben" license="425179">
              <RESULTS>
                <RESULT resultid="1590" eventid="6" swimtime="00:01:30.95" lane="2" heatid="6009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1591" eventid="8" swimtime="00:00:31.59" lane="3" heatid="8019" />
                <RESULT resultid="1592" eventid="10" swimtime="00:01:21.89" lane="2" heatid="10010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="344" birthdate="2015-01-01" gender="F" lastname="Lindner" firstname="Magdalena" license="477898">
              <RESULTS>
                <RESULT resultid="1593" eventid="3" swimtime="00:00:55.52" lane="3" heatid="3004" />
                <RESULT resultid="1594" eventid="7" swimtime="00:00:49.68" lane="1" heatid="7003" />
                <RESULT resultid="1595" eventid="9" swimtime="00:02:14.06" lane="4" heatid="9011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="345" birthdate="2013-01-01" gender="M" lastname="Lindner" firstname="Michael" license="458458">
              <RESULTS>
                <RESULT resultid="1596" eventid="4" swimtime="00:00:48.40" lane="2" heatid="4004" />
                <RESULT resultid="1597" eventid="8" swimtime="00:00:42.57" lane="2" heatid="8005" />
                <RESULT resultid="1598" eventid="10" swimtime="00:01:52.46" lane="1" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="346" birthdate="2011-01-01" gender="F" lastname="Naumann" firstname="Lilly" license="432056">
              <RESULTS>
                <RESULT resultid="1599" eventid="3" swimtime="00:00:44.07" lane="1" heatid="3014" />
                <RESULT resultid="1600" eventid="5" swimtime="00:01:45.06" lane="3" heatid="5006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1601" eventid="9" swimtime="00:01:37.38" lane="2" heatid="9008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="347" birthdate="2011-01-01" gender="F" lastname="Uhlig" firstname="Charlotte" license="446989">
              <RESULTS>
                <RESULT resultid="1602" eventid="5" swimtime="00:01:47.73" lane="2" heatid="5005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1603" eventid="7" swimtime="00:00:45.33" lane="2" heatid="7009" />
                <RESULT resultid="1604" eventid="9" swimtime="00:01:50.21" lane="2" heatid="9005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="348" birthdate="2013-01-01" gender="F" lastname="Uhlig" firstname="Magdalena" license="451879">
              <RESULTS>
                <RESULT resultid="1605" eventid="5" swimtime="00:01:42.47" lane="1" heatid="5010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1606" eventid="7" swimtime="00:00:38.19" lane="4" heatid="7014" />
                <RESULT resultid="1607" eventid="9" swimtime="00:01:35.66" lane="1" heatid="9013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="349" birthdate="2015-01-01" gender="F" lastname="Wendler" firstname="Hilde Ella" license="477900">
              <RESULTS>
                <RESULT resultid="1608" eventid="3" swimtime="00:01:02.24" lane="1" heatid="3002" />
                <RESULT resultid="1609" eventid="5" swimtime="00:02:34.47" lane="1" heatid="5001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1610" eventid="7" swimtime="00:00:59.51" lane="1" heatid="7001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="350" birthdate="2011-01-01" gender="F" lastname="Wolf" firstname="Anastasia" license="425176">
              <RESULTS>
                <RESULT resultid="1611" eventid="3" status="DSQ" swimtime="00:00:43.43" lane="1" heatid="3016" comment="Die Sportlerin hat bei der Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt." />
                <RESULT resultid="1612" eventid="7" swimtime="00:00:35.71" lane="4" heatid="7017" />
                <RESULT resultid="1613" eventid="9" swimtime="00:01:33.05" lane="3" heatid="9009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Weixdorf e.V." nation="GER" region="12" code="3366">
          <ATHLETES>
            <ATHLETE athleteid="40" birthdate="2005-01-01" gender="F" lastname="Conrad" firstname="Linda" license="298857">
              <RESULTS>
                <RESULT resultid="143" eventid="27" swimtime="00:00:36.56" lane="1" heatid="27008" />
                <RESULT resultid="144" eventid="33" swimtime="00:01:12.17" lane="3" heatid="33010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="145" eventid="37" swimtime="00:02:51.24" lane="2" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:21.27" />
                    <SPLIT distance="150" swimtime="00:02:06.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="146" eventid="41" swimtime="00:00:32.55" lane="1" heatid="41008" />
                <RESULT resultid="147" eventid="45" swimtime="00:01:18.86" lane="3" heatid="45006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2059" eventid="60" swimtime="00:00:35.69" lane="1" heatid="60001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="41" birthdate="2004-01-01" gender="F" lastname="Meyer" firstname="Joelle Marie" license="307333">
              <RESULTS>
                <RESULT resultid="148" eventid="25" swimtime="00:00:30.19" lane="2" heatid="25013" />
                <RESULT resultid="149" eventid="29" swimtime="00:01:08.91" lane="2" heatid="29007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="150" eventid="33" swimtime="00:01:09.86" lane="2" heatid="33011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="151" eventid="41" swimtime="00:00:28.67" lane="3" heatid="41014" />
                <RESULT resultid="152" eventid="43" swimtime="00:00:27.65" lane="3" heatid="43017" />
                <RESULT resultid="2043" eventid="56" swimtime="00:00:29.79" lane="1" heatid="56001" />
                <RESULT resultid="2076" eventid="64" swimtime="00:00:28.44" lane="3" heatid="64001" />
                <RESULT resultid="2092" eventid="68" swimtime="00:00:27.65" lane="3" heatid="68001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Würzburg 05" nation="GER" region="2" code="4339">
          <ATHLETES>
            <ATHLETE athleteid="57" birthdate="2009-01-01" gender="M" lastname="Schmidt" firstname="Till Melvin" license="404171">
              <RESULTS>
                <RESULT resultid="228" eventid="30" swimtime="00:01:12.76" lane="4" heatid="30001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="229" eventid="32" swimtime="00:01:02.64" lane="3" heatid="32008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="230" eventid="50" swimtime="00:02:50.34" lane="3" heatid="50001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:19.08" />
                    <SPLIT distance="150" swimtime="00:02:04.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="231" eventid="52" swimtime="00:02:18.01" lane="1" heatid="52004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:06.15" />
                    <SPLIT distance="150" swimtime="00:01:43.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Zwickau von 1904" nation="GER" region="12" code="3400">
          <ATHLETES>
            <ATHLETE athleteid="176" birthdate="2015-01-01" gender="F" lastname="Birzer" firstname="Frieda" license="466284">
              <RESULTS>
                <RESULT resultid="789" eventid="3" swimtime="00:00:48.31" lane="1" heatid="3018" />
                <RESULT resultid="790" eventid="7" swimtime="00:00:44.20" lane="4" heatid="7019" />
                <RESULT resultid="791" eventid="15" swimtime="00:01:46.62" lane="1" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="792" eventid="17" swimtime="00:00:52.71" lane="3" heatid="17010" />
                <RESULT resultid="793" eventid="19" swimtime="00:01:41.00" lane="1" heatid="19003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="177" birthdate="2013-01-01" gender="F" lastname="Dressel" firstname="Clara" license="447504">
              <RESULTS>
                <RESULT resultid="794" eventid="3" swimtime="00:00:44.82" lane="4" heatid="3013" />
                <RESULT resultid="795" eventid="7" swimtime="00:00:38.61" lane="4" heatid="7013" />
                <RESULT resultid="796" eventid="9" swimtime="00:01:37.53" lane="3" heatid="9007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="797" eventid="15" swimtime="00:01:36.27" lane="1" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="798" eventid="19" swimtime="00:01:27.70" lane="4" heatid="19008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="799" eventid="21" swimtime="00:03:29.03" lane="2" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                    <SPLIT distance="100" swimtime="00:01:44.29" />
                    <SPLIT distance="150" swimtime="00:02:44.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="178" birthdate="2015-01-01" gender="F" lastname="Dusl" firstname="Mara" license="466278">
              <RESULTS>
                <RESULT resultid="800" eventid="3" swimtime="00:00:50.40" lane="4" heatid="3006" />
                <RESULT resultid="801" eventid="5" swimtime="00:02:06.65" lane="4" heatid="5008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="802" eventid="15" swimtime="00:01:53.65" lane="4" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="803" eventid="17" swimtime="00:01:00.00" lane="3" heatid="17003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="179" birthdate="2008-01-01" gender="F" lastname="Epperlein" firstname="Linda" license="367581">
              <RESULTS>
                <RESULT resultid="804" eventid="29" status="DNS" swimtime="00:00:00.00" lane="4" heatid="29002" />
                <RESULT resultid="805" eventid="31" status="DNS" swimtime="00:00:00.00" lane="3" heatid="31003" />
                <RESULT resultid="806" eventid="41" status="DNS" swimtime="00:00:00.00" lane="4" heatid="41005" />
                <RESULT resultid="807" eventid="43" status="DNS" swimtime="00:00:00.00" lane="4" heatid="43004" />
                <RESULT resultid="808" eventid="49" status="DNS" swimtime="00:00:00.00" lane="3" heatid="49001" />
                <RESULT resultid="809" eventid="51" status="DNS" swimtime="00:00:00.00" lane="4" heatid="51003" />
                <RESULT resultid="810" eventid="53" status="DNS" swimtime="00:00:00.00" lane="3" heatid="53002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="180" birthdate="2013-01-01" gender="F" lastname="Fenzel" firstname="Valeria" license="448580">
              <RESULTS>
                <RESULT resultid="811" eventid="3" swimtime="00:00:43.47" lane="4" heatid="3014" />
                <RESULT resultid="812" eventid="7" swimtime="00:00:38.08" lane="2" heatid="7014" />
                <RESULT resultid="813" eventid="9" swimtime="00:01:37.63" lane="4" heatid="9013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="814" eventid="13" swimtime="00:00:48.13" lane="4" heatid="13008" />
                <RESULT resultid="815" eventid="15" swimtime="00:01:36.46" lane="4" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="816" eventid="19" swimtime="00:01:28.57" lane="4" heatid="19014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="181" birthdate="2007-01-01" gender="F" lastname="Hupfer" firstname="Louise" license="402573">
              <RESULTS>
                <RESULT resultid="817" eventid="25" status="DNS" swimtime="00:00:00.00" lane="2" heatid="25003" />
                <RESULT resultid="818" eventid="27" status="DNS" swimtime="00:00:00.00" lane="1" heatid="27002" />
                <RESULT resultid="819" eventid="31" status="DNS" swimtime="00:00:00.00" lane="4" heatid="31003" />
                <RESULT resultid="820" eventid="45" status="DNS" swimtime="00:00:00.00" lane="3" heatid="45001" />
                <RESULT resultid="821" eventid="47" status="DNS" swimtime="00:00:00.00" lane="2" heatid="47001" />
                <RESULT resultid="822" eventid="51" status="DNS" swimtime="00:00:00.00" lane="1" heatid="51003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182" birthdate="2003-01-01" gender="F" lastname="Jörg" firstname="Loreen" license="309483">
              <RESULTS>
                <RESULT resultid="823" eventid="27" swimtime="00:00:39.74" lane="3" heatid="27009" />
                <RESULT resultid="824" eventid="29" swimtime="00:01:17.37" lane="3" heatid="29002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="825" eventid="31" swimtime="00:01:10.95" lane="3" heatid="31007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="826" eventid="41" swimtime="00:00:33.86" lane="2" heatid="41008" />
                <RESULT resultid="827" eventid="43" swimtime="00:00:31.70" lane="4" heatid="43008" />
                <RESULT resultid="828" eventid="45" swimtime="00:01:25.95" lane="3" heatid="45007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183" birthdate="2010-01-01" gender="M" lastname="Käser" firstname="Mika Marco" license="423052">
              <RESULTS>
                <RESULT resultid="829" eventid="6" swimtime="00:01:30.55" lane="3" heatid="6010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="830" eventid="8" swimtime="00:00:31.44" lane="2" heatid="8014" />
                <RESULT resultid="831" eventid="10" swimtime="00:01:22.27" lane="4" heatid="10011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="832" eventid="16" swimtime="00:01:21.41" lane="3" heatid="16009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="833" eventid="18" swimtime="00:00:42.22" lane="1" heatid="18013" />
                <RESULT resultid="834" eventid="20" swimtime="00:01:12.35" lane="4" heatid="20016">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="184" birthdate="2007-01-01" gender="F" lastname="Klose" firstname="Klara" license="364236">
              <RESULTS>
                <RESULT resultid="835" eventid="25" swimtime="00:00:38.30" lane="1" heatid="25005" />
                <RESULT resultid="836" eventid="27" swimtime="00:00:42.57" lane="3" heatid="27003" />
                <RESULT resultid="837" eventid="31" swimtime="00:01:12.33" lane="1" heatid="31006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="838" eventid="43" swimtime="00:00:31.19" lane="2" heatid="43010" />
                <RESULT resultid="839" eventid="47" swimtime="00:01:26.70" lane="2" heatid="47004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="185" birthdate="2012-01-01" gender="F" lastname="Komar" firstname="Lindsay" license="436924">
              <RESULTS>
                <RESULT resultid="840" eventid="1" swimtime="00:01:28.12" lane="4" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="841" eventid="7" swimtime="00:00:34.21" lane="2" heatid="7017" />
                <RESULT resultid="842" eventid="9" swimtime="00:01:26.93" lane="1" heatid="9010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="843" eventid="13" swimtime="00:00:37.02" lane="3" heatid="13009" />
                <RESULT resultid="844" eventid="19" swimtime="00:01:18.63" lane="4" heatid="19011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="845" eventid="21" swimtime="00:03:07.15" lane="4" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:01:27.02" />
                    <SPLIT distance="150" swimtime="00:02:23.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="186" birthdate="2007-01-01" gender="F" lastname="Kunz" firstname="Jenny" license="363787">
              <RESULTS>
                <RESULT resultid="846" eventid="29" status="DNS" swimtime="00:00:00.00" lane="1" heatid="29005" />
                <RESULT resultid="847" eventid="31" status="DNS" swimtime="00:00:00.00" lane="2" heatid="31007" />
                <RESULT resultid="848" eventid="33" status="DNS" swimtime="00:00:00.00" lane="3" heatid="33009" />
                <RESULT resultid="849" eventid="41" status="DNS" swimtime="00:00:00.00" lane="1" heatid="41009" />
                <RESULT resultid="850" eventid="53" status="DNS" swimtime="00:00:00.00" lane="2" heatid="53004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="187" birthdate="2005-01-01" gender="M" lastname="Kunz" firstname="Jeremy" license="348770">
              <RESULTS>
                <RESULT resultid="851" eventid="26" swimtime="00:00:27.62" lane="2" heatid="26010" />
                <RESULT resultid="852" eventid="28" swimtime="00:00:30.85" lane="3" heatid="28008" />
                <RESULT resultid="853" eventid="34" swimtime="00:00:59.35" lane="2" heatid="34007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="854" eventid="42" swimtime="00:00:26.80" lane="4" heatid="42011" />
                <RESULT resultid="855" eventid="44" swimtime="00:00:25.20" lane="2" heatid="44010" />
                <RESULT resultid="856" eventid="52" swimtime="00:01:58.19" lane="2" heatid="52005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="100" swimtime="00:00:59.10" />
                    <SPLIT distance="150" swimtime="00:01:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="857" eventid="54" swimtime="00:02:18.11" lane="2" heatid="54003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2051" eventid="58" swimtime="00:00:27.98" lane="1" heatid="58001" />
                <RESULT resultid="2069" eventid="62" swimtime="00:00:30.97" lane="1" heatid="62001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="188" birthdate="2015-01-01" gender="F" lastname="Lemke" firstname="Lilly-Rose" license="466280">
              <RESULTS>
                <RESULT resultid="858" eventid="3" swimtime="00:00:55.01" lane="4" heatid="3018" />
                <RESULT resultid="859" eventid="7" swimtime="00:00:49.10" lane="4" heatid="7004" />
                <RESULT resultid="860" eventid="17" swimtime="00:01:04.72" lane="1" heatid="17003" />
                <RESULT resultid="861" eventid="19" swimtime="00:02:01.76" lane="1" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="189" birthdate="2000-01-01" gender="F" lastname="Massier" firstname="Vivienne" license="295584">
              <RESULTS>
                <RESULT resultid="862" eventid="27" swimtime="00:00:41.64" lane="4" heatid="27009" />
                <RESULT resultid="863" eventid="31" swimtime="00:01:13.34" lane="4" heatid="31006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="864" eventid="43" swimtime="00:00:31.98" lane="1" heatid="43008" />
                <RESULT resultid="865" eventid="45" swimtime="00:01:35.70" lane="1" heatid="45007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="190" birthdate="2014-01-01" gender="F" lastname="Mittenzwei" firstname="Charlotta" license="456274">
              <RESULTS>
                <RESULT resultid="866" eventid="5" status="DSQ" swimtime="00:01:50.30" lane="3" heatid="5009" comment="Die Sportlerin startete vor dem Startsignal">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="867" eventid="7" swimtime="00:00:43.08" lane="3" heatid="7009" />
                <RESULT resultid="868" eventid="9" swimtime="00:01:49.58" lane="3" heatid="9005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="869" eventid="13" swimtime="00:00:56.13" lane="4" heatid="13007" />
                <RESULT resultid="870" eventid="17" swimtime="00:00:52.14" lane="3" heatid="17011" />
                <RESULT resultid="871" eventid="19" swimtime="00:01:39.37" lane="2" heatid="19004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191" birthdate="2009-01-01" gender="F" lastname="Nahlovsky" firstname="Lilly" license="410485">
              <RESULTS>
                <RESULT resultid="872" eventid="25" swimtime="00:00:31.61" lane="3" heatid="25010" />
                <RESULT resultid="873" eventid="27" swimtime="00:00:38.15" lane="3" heatid="27006" />
                <RESULT resultid="874" eventid="31" swimtime="00:01:04.59" lane="1" heatid="31010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="875" eventid="33" swimtime="00:01:11.63" lane="2" heatid="33008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="876" eventid="41" swimtime="00:00:32.17" lane="1" heatid="41011" />
                <RESULT resultid="877" eventid="43" swimtime="00:00:28.65" lane="2" heatid="43014" />
                <RESULT resultid="878" eventid="47" swimtime="00:01:10.01" lane="3" heatid="47007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2038" eventid="55" swimtime="00:00:31.62" lane="3" heatid="55001" />
                <RESULT resultid="2055" eventid="59" swimtime="00:00:38.00" lane="1" heatid="59001" />
                <RESULT resultid="2089" eventid="67" swimtime="00:00:28.62" lane="1" heatid="67001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="192" birthdate="2012-01-01" gender="M" lastname="Nawrath" firstname="Jonas" license="443627">
              <RESULTS>
                <RESULT resultid="879" eventid="6" swimtime="00:01:39.26" lane="2" heatid="6005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="880" eventid="8" swimtime="00:00:36.37" lane="1" heatid="8010" />
                <RESULT resultid="881" eventid="14" swimtime="00:00:44.40" lane="4" heatid="14006" />
                <RESULT resultid="882" eventid="18" swimtime="00:00:43.36" lane="4" heatid="18011" />
                <RESULT resultid="883" eventid="20" swimtime="00:01:22.13" lane="2" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="884" eventid="22" status="DSQ" swimtime="00:03:19.70" lane="2" heatid="22001" comment="Der Sportler war beim Zielanschlag der Teilstrecke Rücken nicht in Rückenlage.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:36.39" />
                    <SPLIT distance="150" swimtime="00:02:32.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="193" birthdate="2013-01-01" gender="M" lastname="Opitz" firstname="Theodor" license="461990">
              <RESULTS>
                <RESULT resultid="885" eventid="4" swimtime="00:00:49.68" lane="3" heatid="4004" />
                <RESULT resultid="886" eventid="8" swimtime="00:00:48.07" lane="3" heatid="8001" />
                <RESULT resultid="887" eventid="18" swimtime="00:00:53.03" lane="3" heatid="18004" />
                <RESULT resultid="888" eventid="20" swimtime="00:01:59.68" lane="3" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="194" birthdate="2009-01-01" gender="M" lastname="Parthier" firstname="Louis" license="410488">
              <RESULTS>
                <RESULT resultid="889" eventid="26" swimtime="00:00:35.38" lane="1" heatid="26003" />
                <RESULT resultid="890" eventid="32" swimtime="00:01:11.80" lane="4" heatid="32002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="891" eventid="36" swimtime="00:02:46.35" lane="3" heatid="36001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:01:24.59" />
                    <SPLIT distance="150" swimtime="00:02:07.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="892" eventid="44" swimtime="00:00:31.71" lane="2" heatid="44001" />
                <RESULT resultid="893" eventid="48" swimtime="00:01:16.83" lane="1" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195" birthdate="2004-01-01" gender="M" lastname="Paul" firstname="Lenny" license="331135">
              <RESULTS>
                <RESULT resultid="894" eventid="26" swimtime="00:00:30.70" lane="2" heatid="26005" />
                <RESULT resultid="895" eventid="28" swimtime="00:00:34.15" lane="4" heatid="28005" />
                <RESULT resultid="896" eventid="30" swimtime="00:01:02.49" lane="4" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="897" eventid="34" swimtime="00:01:07.86" lane="2" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="898" eventid="42" swimtime="00:00:27.58" lane="3" heatid="42008" />
                <RESULT resultid="899" eventid="46" swimtime="00:01:18.19" lane="1" heatid="46006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196" birthdate="2003-01-01" gender="F" lastname="Pelloth" firstname="Anne-Katrin" license="365577">
              <RESULTS>
                <RESULT resultid="900" eventid="25" swimtime="00:00:34.71" lane="3" heatid="25007" />
                <RESULT resultid="901" eventid="29" swimtime="00:01:14.09" lane="1" heatid="29007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="902" eventid="31" swimtime="00:01:05.61" lane="2" heatid="31013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="903" eventid="33" swimtime="00:01:15.95" lane="3" heatid="33011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="904" eventid="41" swimtime="00:00:32.63" lane="4" heatid="41014" />
                <RESULT resultid="905" eventid="43" swimtime="00:00:29.59" lane="4" heatid="43017" />
                <RESULT resultid="906" eventid="53" swimtime="00:02:46.75" lane="3" heatid="53004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:15.48" />
                    <SPLIT distance="150" swimtime="00:02:05.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197" birthdate="2014-01-01" gender="M" lastname="Plettig" firstname="Ben" license="464151">
              <RESULTS>
                <RESULT resultid="907" eventid="4" swimtime="00:00:46.88" lane="4" heatid="4011" />
                <RESULT resultid="908" eventid="8" swimtime="00:00:44.05" lane="1" heatid="8005" />
                <RESULT resultid="909" eventid="10" swimtime="00:01:47.85" lane="3" heatid="10007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="910" eventid="18" swimtime="00:00:59.49" lane="3" heatid="18002" />
                <RESULT resultid="911" eventid="20" swimtime="00:01:37.40" lane="2" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198" birthdate="2006-01-01" gender="F" lastname="Rebentisch" firstname="Maya" license="342540">
              <RESULTS>
                <RESULT resultid="912" eventid="25" swimtime="00:00:39.15" lane="4" heatid="25012" />
                <RESULT resultid="913" eventid="33" swimtime="00:01:35.61" lane="4" heatid="33010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="914" eventid="35" swimtime="00:03:07.42" lane="2" heatid="35001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                    <SPLIT distance="100" swimtime="00:01:32.97" />
                    <SPLIT distance="150" swimtime="00:02:22.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="915" eventid="43" swimtime="00:00:37.50" lane="4" heatid="43002" />
                <RESULT resultid="916" eventid="47" status="DSQ" swimtime="00:01:26.99" lane="1" heatid="47009" comment="Die Sportlerin hat bei der zweiten Wende nach Verlassen der Rückenlage nicht unverzüglich die eigentliche Wendenbewegung ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="199" birthdate="2013-01-01" gender="M" lastname="Richter" firstname="Luke" license="446150">
              <RESULTS>
                <RESULT resultid="917" eventid="4" swimtime="00:00:41.66" lane="4" heatid="4012" />
                <RESULT resultid="918" eventid="8" swimtime="00:00:34.87" lane="1" heatid="8017" />
                <RESULT resultid="919" eventid="10" swimtime="00:01:35.55" lane="4" heatid="10005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="920" eventid="14" status="DNS" swimtime="00:00:00.00" lane="1" heatid="14005" />
                <RESULT resultid="921" eventid="16" swimtime="00:01:32.09" lane="2" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="922" eventid="20" swimtime="00:01:23.01" lane="4" heatid="20010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="200" birthdate="2010-01-01" gender="F" lastname="Rohatzsch" firstname="Maxime" license="410491">
              <RESULTS>
                <RESULT resultid="923" eventid="25" swimtime="00:00:35.11" lane="1" heatid="25009" />
                <RESULT resultid="924" eventid="29" swimtime="00:01:29.75" lane="1" heatid="29003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="925" eventid="33" swimtime="00:01:19.05" lane="1" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="926" eventid="35" swimtime="00:02:49.44" lane="3" heatid="35002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:21.25" />
                    <SPLIT distance="150" swimtime="00:02:06.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="927" eventid="41" swimtime="00:00:37.48" lane="3" heatid="41010" />
                <RESULT resultid="928" eventid="47" swimtime="00:01:18.44" lane="3" heatid="47006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="929" eventid="53" status="DNS" swimtime="00:00:00.00" lane="2" heatid="53003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201" birthdate="1999-01-01" gender="M" lastname="Schneider" firstname="Eric" license="242941">
              <RESULTS>
                <RESULT resultid="930" eventid="26" swimtime="00:00:28.21" lane="3" heatid="26007" />
                <RESULT resultid="931" eventid="28" swimtime="00:00:31.71" lane="1" heatid="28009" />
                <RESULT resultid="932" eventid="34" swimtime="00:01:01.22" lane="3" heatid="34008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="933" eventid="42" swimtime="00:00:26.94" lane="2" heatid="42008" />
                <RESULT resultid="934" eventid="44" swimtime="00:00:25.26" lane="3" heatid="44010" />
                <RESULT resultid="2052" eventid="58" swimtime="00:00:28.35" lane="4" heatid="58001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202" birthdate="2013-01-01" gender="F" lastname="Schneider" firstname="Laura" license="447503">
              <RESULTS>
                <RESULT resultid="935" eventid="3" swimtime="00:00:39.01" lane="2" heatid="3020" />
                <RESULT resultid="936" eventid="5" swimtime="00:01:35.53" lane="2" heatid="5010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="937" eventid="9" swimtime="00:01:29.36" lane="3" heatid="9013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="938" eventid="13" status="DNS" swimtime="00:00:00.00" lane="2" heatid="13008" />
                <RESULT resultid="939" eventid="17" swimtime="00:00:42.88" lane="2" heatid="17012" />
                <RESULT resultid="940" eventid="21" swimtime="00:03:12.93" lane="2" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                    <SPLIT distance="100" swimtime="00:01:31.77" />
                    <SPLIT distance="150" swimtime="00:02:27.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="203" birthdate="2007-01-01" gender="F" lastname="Schneider" firstname="Shanya" license="394943">
              <RESULTS>
                <RESULT resultid="941" eventid="25" swimtime="00:00:39.20" lane="2" heatid="25004" />
                <RESULT resultid="942" eventid="27" swimtime="00:00:44.11" lane="1" heatid="27003" />
                <RESULT resultid="943" eventid="31" swimtime="00:01:17.69" lane="2" heatid="31003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="944" eventid="33" swimtime="00:01:25.08" lane="3" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="945" eventid="41" swimtime="00:00:36.81" lane="2" heatid="41004" />
                <RESULT resultid="946" eventid="43" swimtime="00:00:33.97" lane="2" heatid="43005" />
                <RESULT resultid="947" eventid="47" swimtime="00:01:25.24" lane="2" heatid="47003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="204" birthdate="2009-01-01" gender="M" lastname="Schulz" firstname="Laurenz" license="394944">
              <RESULTS>
                <RESULT resultid="948" eventid="26" swimtime="00:00:33.12" lane="3" heatid="26008" />
                <RESULT resultid="949" eventid="30" swimtime="00:01:14.37" lane="2" heatid="30001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="950" eventid="34" swimtime="00:01:17.86" lane="3" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="951" eventid="42" swimtime="00:00:31.51" lane="3" heatid="42009" />
                <RESULT resultid="952" eventid="48" swimtime="00:01:16.51" lane="3" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="953" eventid="54" swimtime="00:02:46.74" lane="2" heatid="54001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                    <SPLIT distance="150" swimtime="00:02:07.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="205" birthdate="2014-01-01" gender="F" lastname="Sprenger" firstname="Lara" license="456271">
              <RESULTS>
                <RESULT resultid="954" eventid="3" swimtime="00:00:45.74" lane="1" heatid="3019" />
                <RESULT resultid="955" eventid="7" swimtime="00:00:40.09" lane="1" heatid="7020" />
                <RESULT resultid="956" eventid="9" swimtime="00:01:48.13" lane="4" heatid="9012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="957" eventid="13" swimtime="00:00:54.33" lane="2" heatid="13001" />
                <RESULT resultid="958" eventid="15" swimtime="00:01:45.11" lane="1" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="959" eventid="19" swimtime="00:01:41.13" lane="1" heatid="19013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="206" birthdate="2010-01-01" gender="M" lastname="Sprenger" firstname="Tom" license="416252">
              <RESULTS>
                <RESULT resultid="960" eventid="4" swimtime="00:00:42.66" lane="1" heatid="4008" />
                <RESULT resultid="961" eventid="8" swimtime="00:00:35.36" lane="4" heatid="8013" />
                <RESULT resultid="962" eventid="10" status="DSQ" swimtime="00:01:35.23" lane="1" heatid="10005" comment="Auf der Teilstrecke Brust wurden die Füße in der Rückwärtsbewegung des beinschlags nicht auswärts gedreht.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="963" eventid="16" swimtime="00:01:34.81" lane="4" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="964" eventid="20" swimtime="00:01:18.52" lane="2" heatid="20009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="207" birthdate="2004-01-01" gender="F" lastname="Süppel" firstname="Laura" license="329276">
              <RESULTS>
                <RESULT resultid="965" eventid="25" swimtime="00:00:35.82" lane="3" heatid="25006" />
                <RESULT resultid="966" eventid="29" swimtime="00:01:18.43" lane="4" heatid="29007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="967" eventid="31" swimtime="00:01:13.77" lane="4" heatid="31007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="968" eventid="33" swimtime="00:01:18.97" lane="4" heatid="33011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="969" eventid="41" swimtime="00:00:32.80" lane="4" heatid="41009" />
                <RESULT resultid="970" eventid="47" swimtime="00:01:18.95" lane="4" heatid="47010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="971" eventid="53" swimtime="00:02:52.45" lane="4" heatid="53004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                    <SPLIT distance="150" swimtime="00:02:11.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="208" birthdate="2004-01-01" gender="M" lastname="Walther" firstname="Theo" license="314090">
              <RESULTS>
                <RESULT resultid="972" eventid="26" swimtime="00:00:29.86" lane="1" heatid="26006" />
                <RESULT resultid="973" eventid="32" swimtime="00:00:59.54" lane="1" heatid="32011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="974" eventid="42" swimtime="00:00:29.69" lane="3" heatid="42006" />
                <RESULT resultid="975" eventid="44" swimtime="00:00:27.59" lane="4" heatid="44008" />
                <RESULT resultid="976" eventid="46" swimtime="00:01:19.43" lane="4" heatid="46006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="977" eventid="48" swimtime="00:01:09.14" lane="4" heatid="48006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="209" birthdate="2011-01-01" gender="M" lastname="Wölki" firstname="Luca" license="430687">
              <RESULTS>
                <RESULT resultid="978" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="979" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="980" eventid="10" status="WDR" swimtime="00:00:00.00" lane="0" heatid="10000" />
                <RESULT resultid="981" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="982" eventid="18" status="WDR" swimtime="00:00:00.00" lane="0" heatid="18000" />
                <RESULT resultid="983" eventid="20" status="WDR" swimtime="00:00:00.00" lane="0" heatid="20000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210" birthdate="2013-01-01" gender="F" lastname="Zaiaieva" firstname="Vlada" license="468008">
              <RESULTS>
                <RESULT resultid="984" eventid="3" swimtime="00:00:47.40" lane="2" heatid="3012" />
                <RESULT resultid="985" eventid="7" swimtime="00:00:40.50" lane="1" heatid="7012" />
                <RESULT resultid="986" eventid="9" status="DSQ" swimtime="00:01:47.95" lane="1" heatid="9007" comment="Die Sportlerin hat die Teilstrecke Rücken nicht in Rückenlage.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="987" eventid="15" swimtime="00:01:42.24" lane="3" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="988" eventid="17" swimtime="00:00:58.55" lane="2" heatid="17003" />
                <RESULT resultid="989" eventid="19" swimtime="00:01:32.06" lane="2" heatid="19007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="211" birthdate="2014-01-01" gender="M" lastname="Zänsler" firstname="Elias" license="461989">
              <RESULTS>
                <RESULT resultid="990" eventid="4" swimtime="00:00:51.23" lane="2" heatid="4002" />
                <RESULT resultid="991" eventid="8" swimtime="00:03:49.60" lane="3" heatid="8004" />
                <RESULT resultid="992" eventid="10" swimtime="00:01:57.08" lane="4" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="993" eventid="20" swimtime="00:01:57.88" lane="4" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="783" eventid="40" swimtime="00:01:41.82" lane="1" heatid="40003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="100" swimtime="00:00:51.47" />
                    <SPLIT distance="150" swimtime="00:01:17.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="208" number="1" />
                    <RELAYPOSITION athleteid="201" number="2" />
                    <RELAYPOSITION athleteid="195" number="3" />
                    <RELAYPOSITION athleteid="187" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="784" eventid="72" swimtime="00:01:51.03" lane="1" heatid="72003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="100" swimtime="00:00:59.42" />
                    <SPLIT distance="150" swimtime="00:01:26.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="208" number="1" />
                    <RELAYPOSITION athleteid="187" number="2" />
                    <RELAYPOSITION athleteid="195" number="3" />
                    <RELAYPOSITION athleteid="201" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="785" eventid="39" swimtime="00:01:59.53" lane="2" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:01:00.27" />
                    <SPLIT distance="150" swimtime="00:01:31.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="196" number="1" />
                    <RELAYPOSITION athleteid="184" number="2" />
                    <RELAYPOSITION athleteid="182" number="3" />
                    <RELAYPOSITION athleteid="191" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="786" eventid="71" swimtime="00:02:13.53" lane="1" heatid="71003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                    <SPLIT distance="150" swimtime="00:01:45.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="196" number="1" />
                    <RELAYPOSITION athleteid="182" number="2" />
                    <RELAYPOSITION athleteid="207" number="3" />
                    <RELAYPOSITION athleteid="191" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="787" eventid="11" swimtime="00:02:11.83" lane="2" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:06.90" />
                    <SPLIT distance="150" swimtime="00:01:40.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="200" number="1" />
                    <RELAYPOSITION athleteid="199" number="2" />
                    <RELAYPOSITION athleteid="185" number="3" />
                    <RELAYPOSITION athleteid="183" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="788" eventid="23" swimtime="00:02:28.58" lane="3" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:22.73" />
                    <SPLIT distance="150" swimtime="00:01:58.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="185" number="1" />
                    <RELAYPOSITION athleteid="202" number="2" />
                    <RELAYPOSITION athleteid="200" number="3" />
                    <RELAYPOSITION athleteid="183" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SV07 Annaberg-Buchholz" nation="GER" region="12" code="3380">
          <ATHLETES>
            <ATHLETE athleteid="321" birthdate="2006-01-01" gender="M" lastname="Schauer" firstname="Lukas" license="365572">
              <RESULTS>
                <RESULT resultid="1478" eventid="26" swimtime="00:00:31.95" lane="3" heatid="26005" />
                <RESULT resultid="1479" eventid="34" swimtime="00:01:12.07" lane="1" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1480" eventid="42" swimtime="00:00:29.48" lane="1" heatid="42005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="322" birthdate="2005-01-01" gender="M" lastname="Siegel" firstname="Paul" license="343558">
              <RESULTS>
                <RESULT resultid="1481" eventid="26" swimtime="00:00:31.63" lane="4" heatid="26005" />
                <RESULT resultid="1482" eventid="32" swimtime="00:00:55.93" lane="2" heatid="32007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1483" eventid="44" swimtime="00:00:25.25" lane="3" heatid="44013" />
                <RESULT resultid="1484" eventid="48" swimtime="00:01:10.59" lane="4" heatid="48005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SVV Plauen" nation="GER" region="12" code="6253">
          <ATHLETES>
            <ATHLETE athleteid="2" birthdate="2012-01-01" gender="M" lastname="Lindner" firstname="Laurence" license="439928">
              <RESULTS>
                <RESULT resultid="8" eventid="2" swimtime="00:01:15.21" lane="2" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="9" eventid="10" swimtime="00:01:16.53" lane="3" heatid="10009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="10" eventid="14" swimtime="00:00:33.99" lane="2" heatid="14009" />
                <RESULT resultid="11" eventid="22" status="DNS" swimtime="00:00:00.00" lane="2" heatid="22003" />
                <RESULT resultid="12" eventid="36" status="DNS" swimtime="00:00:00.00" lane="2" heatid="36001" />
                <RESULT resultid="13" eventid="52" status="DNS" swimtime="00:00:00.00" lane="3" heatid="52003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="3" birthdate="2012-01-01" gender="M" lastname="Mocker" firstname="Felix" license="439927">
              <RESULTS>
                <RESULT resultid="14" eventid="6" swimtime="00:01:27.76" lane="3" heatid="6008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="15" eventid="10" swimtime="00:01:21.19" lane="4" heatid="10009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="16" eventid="16" swimtime="00:01:23.60" lane="2" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="17" eventid="18" swimtime="00:00:42.00" lane="3" heatid="18011" />
                <RESULT resultid="18" eventid="38" swimtime="00:03:05.79" lane="1" heatid="38001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:29.22" />
                    <SPLIT distance="150" swimtime="00:02:17.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="19" eventid="52" swimtime="00:02:36.96" lane="1" heatid="52002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:57.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TJ Slavie Chomutov" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="266" birthdate="2007-01-01" gender="F" lastname="Doksanská" firstname="Anezka" license="0">
              <RESULTS>
                <RESULT resultid="1203" eventid="25" swimtime="00:00:31.44" lane="2" heatid="25011" />
                <RESULT resultid="1204" eventid="31" swimtime="00:01:03.52" lane="4" heatid="31011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1205" eventid="35" swimtime="00:02:26.87" lane="2" heatid="35003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:50.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1206" eventid="43" swimtime="00:00:28.95" lane="4" heatid="43015" />
                <RESULT resultid="1207" eventid="47" swimtime="00:01:07.50" lane="2" heatid="47008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2037" eventid="55" swimtime="00:00:31.18" lane="2" heatid="55001" />
                <RESULT resultid="2090" eventid="67" swimtime="00:00:28.61" lane="4" heatid="67001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="267" birthdate="2008-01-01" gender="F" lastname="Hájková" firstname="Marie" license="0">
              <RESULTS>
                <RESULT resultid="1209" eventid="27" status="DNS" swimtime="00:00:00.00" lane="4" heatid="27002" />
                <RESULT resultid="1210" eventid="31" swimtime="00:01:16.20" lane="1" heatid="31007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1212" eventid="33" swimtime="00:01:30.82" lane="4" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1211" eventid="43" swimtime="00:00:34.81" lane="4" heatid="43009" />
                <RESULT resultid="1213" eventid="45" status="DNS" swimtime="00:00:00.00" lane="2" heatid="45001" />
                <RESULT resultid="1208" eventid="47" swimtime="00:01:34.99" lane="3" heatid="47004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="268" birthdate="2008-01-01" gender="F" lastname="Jirová" firstname="Petra" license="0">
              <RESULTS>
                <RESULT resultid="1214" eventid="25" status="DNS" swimtime="00:00:00.00" lane="2" heatid="25006" />
                <RESULT resultid="1215" eventid="31" status="DNS" swimtime="00:00:00.00" lane="2" heatid="31008" />
                <RESULT resultid="1216" eventid="33" status="DNS" swimtime="00:00:00.00" lane="2" heatid="33009" />
                <RESULT resultid="1217" eventid="41" status="DNS" swimtime="00:00:00.00" lane="1" heatid="41012" />
                <RESULT resultid="1218" eventid="43" status="DNS" swimtime="00:00:00.00" lane="1" heatid="43012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="269" birthdate="2002-01-01" gender="F" lastname="Malinová" firstname="Michaela" license="0">
              <RESULTS>
                <RESULT resultid="1219" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="1220" eventid="33" status="WDR" swimtime="00:00:00.00" lane="0" heatid="33000" />
                <RESULT resultid="1221" eventid="43" status="WDR" swimtime="00:00:00.00" lane="0" heatid="43000" />
                <RESULT resultid="1222" eventid="45" status="WDR" swimtime="00:00:00.00" lane="0" heatid="45000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="270" birthdate="2007-01-01" gender="F" lastname="Nevolová" firstname="Katerina" license="0">
              <RESULTS>
                <RESULT resultid="1223" eventid="25" swimtime="00:00:33.38" lane="1" heatid="25008" />
                <RESULT resultid="1224" eventid="31" swimtime="00:01:05.86" lane="3" heatid="31008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1225" eventid="35" swimtime="00:02:33.64" lane="1" heatid="35003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="150" swimtime="00:01:54.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1226" eventid="43" swimtime="00:00:30.25" lane="4" heatid="43011" />
                <RESULT resultid="1227" eventid="47" swimtime="00:01:11.08" lane="1" heatid="47008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="271" birthdate="2005-01-01" gender="F" lastname="Svobodová" firstname="Zuzana" license="0">
              <RESULTS>
                <RESULT resultid="1228" eventid="27" swimtime="00:00:34.84" lane="3" heatid="27008" />
                <RESULT resultid="1229" eventid="33" swimtime="00:01:13.69" lane="2" heatid="33010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1230" eventid="37" swimtime="00:02:51.98" lane="3" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:01:22.98" />
                    <SPLIT distance="150" swimtime="00:02:08.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1231" eventid="41" swimtime="00:00:34.60" lane="2" heatid="41005" />
                <RESULT resultid="1232" eventid="43" swimtime="00:00:29.97" lane="1" heatid="43016" />
                <RESULT resultid="1233" eventid="45" swimtime="00:01:18.08" lane="2" heatid="45006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1234" eventid="53" status="DNS" swimtime="00:00:00.00" lane="4" heatid="53005" />
                <RESULT resultid="2057" eventid="60" swimtime="00:00:34.68" lane="2" heatid="60001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="272" birthdate="2008-01-01" gender="F" lastname="Tautrmanová" firstname="Katerina" license="0">
              <RESULTS>
                <RESULT resultid="1235" eventid="25" swimtime="00:00:32.57" lane="2" heatid="25008" />
                <RESULT resultid="1236" eventid="31" swimtime="00:01:01.80" lane="3" heatid="31011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1237" eventid="43" swimtime="00:00:27.94" lane="2" heatid="43015" />
                <RESULT resultid="1238" eventid="47" swimtime="00:01:09.70" lane="3" heatid="47008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1239" eventid="51" swimtime="00:02:15.74" lane="2" heatid="51005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="100" swimtime="00:01:05.38" />
                    <SPLIT distance="150" swimtime="00:01:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2087" eventid="67" swimtime="00:00:27.67" lane="2" heatid="67001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="273" birthdate="2007-01-01" gender="F" lastname="Vlasáková" firstname="Tereza" license="0">
              <RESULTS>
                <RESULT resultid="1240" eventid="25" swimtime="00:00:32.55" lane="4" heatid="25011" />
                <RESULT resultid="1241" eventid="29" status="DNS" swimtime="00:00:00.00" lane="2" heatid="29005" />
                <RESULT resultid="1242" eventid="31" status="DNS" swimtime="00:00:00.00" lane="1" heatid="31011" />
                <RESULT resultid="1243" eventid="41" swimtime="00:00:30.28" lane="2" heatid="41012" />
                <RESULT resultid="1244" eventid="49" swimtime="00:02:33.64" lane="3" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="150" swimtime="00:01:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1245" eventid="53" swimtime="00:02:36.21" lane="3" heatid="53005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:14.52" />
                    <SPLIT distance="150" swimtime="00:01:59.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2040" eventid="55" swimtime="00:00:32.47" lane="4" heatid="55001" />
                <RESULT resultid="2071" eventid="63" swimtime="00:00:30.27" lane="2" heatid="63001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="274" birthdate="2010-01-01" gender="F" lastname="Hájková" firstname="Katerina" license="0">
              <RESULTS>
                <RESULT resultid="1246" eventid="29" swimtime="00:01:38.98" lane="1" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1247" eventid="31" swimtime="00:01:20.19" lane="1" heatid="31009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1248" eventid="33" swimtime="00:01:30.57" lane="2" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1249" eventid="41" swimtime="00:00:42.21" lane="3" heatid="41003" />
                <RESULT resultid="1250" eventid="43" swimtime="00:00:36.05" lane="1" heatid="43004" />
                <RESULT resultid="1251" eventid="49" swimtime="00:03:51.86" lane="1" heatid="49001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:38.81" />
                    <SPLIT distance="150" swimtime="00:02:44.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="275" birthdate="2002-01-01" gender="M" lastname="Jezbera" firstname="Filip" license="0">
              <RESULTS>
                <RESULT resultid="1252" eventid="26" status="WDR" swimtime="00:00:00.00" lane="0" heatid="26000" />
                <RESULT resultid="1253" eventid="44" status="WDR" swimtime="00:00:00.00" lane="0" heatid="44000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="276" birthdate="2007-01-01" gender="M" lastname="Jezbera" firstname="Jakub" license="0">
              <RESULTS>
                <RESULT resultid="1254" eventid="26" swimtime="00:00:30.77" lane="4" heatid="26009" />
                <RESULT resultid="1255" eventid="30" swimtime="00:01:06.10" lane="4" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1256" eventid="32" swimtime="00:01:00.95" lane="4" heatid="32004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1257" eventid="42" swimtime="00:00:30.32" lane="3" heatid="42005" />
                <RESULT resultid="1939" eventid="48" swimtime="00:01:04.71" lane="3" heatid="48004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="277" birthdate="2003-01-01" gender="M" lastname="Kaska" firstname="Karel" license="0">
              <RESULTS>
                <RESULT resultid="1259" eventid="26" swimtime="00:00:28.73" lane="1" heatid="26011" />
                <RESULT resultid="1260" eventid="34" swimtime="00:01:07.78" lane="2" heatid="34008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1261" eventid="44" swimtime="00:00:27.49" lane="3" heatid="44009" />
                <RESULT resultid="1262" eventid="48" swimtime="00:01:03.48" lane="2" heatid="48006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="278" birthdate="2008-01-01" gender="M" lastname="Kubista" firstname="Jan" license="0">
              <RESULTS>
                <RESULT resultid="1263" eventid="26" swimtime="00:00:28.32" lane="2" heatid="26009" />
                <RESULT resultid="1264" eventid="28" swimtime="00:00:33.42" lane="3" heatid="28007" />
                <RESULT resultid="1265" eventid="34" swimtime="00:01:05.73" lane="2" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1266" eventid="44" swimtime="00:00:24.17" lane="2" heatid="44012" />
                <RESULT resultid="1267" eventid="48" swimtime="00:01:05.64" lane="2" heatid="48004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2045" eventid="57" swimtime="00:00:27.19" lane="2" heatid="57001" />
                <RESULT resultid="2063" eventid="61" swimtime="00:00:32.71" lane="3" heatid="61001" />
                <RESULT resultid="2102" eventid="70" swimtime="00:00:24.48" lane="1" heatid="70001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="279" birthdate="2005-01-01" gender="M" lastname="Moravec" firstname="Tomás" license="0">
              <RESULTS>
                <RESULT resultid="1268" eventid="26" swimtime="00:00:28.93" lane="4" heatid="26010" />
                <RESULT resultid="1269" eventid="28" swimtime="00:00:30.40" lane="2" heatid="28008" />
                <RESULT resultid="1270" eventid="32" swimtime="00:00:55.58" lane="2" heatid="32010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1271" eventid="38" swimtime="00:02:21.03" lane="2" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:07.01" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1272" eventid="42" swimtime="00:00:29.83" lane="1" heatid="42008" />
                <RESULT resultid="1273" eventid="46" swimtime="00:01:06.12" lane="2" heatid="46005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2068" eventid="62" swimtime="00:00:30.08" lane="3" heatid="62001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="280" birthdate="2009-01-01" gender="M" lastname="Ocásek" firstname="Daniel" license="0">
              <RESULTS>
                <RESULT resultid="1274" eventid="26" swimtime="00:00:37.88" lane="1" heatid="26001" />
                <RESULT resultid="1275" eventid="28" swimtime="00:00:45.71" lane="3" heatid="28001" />
                <RESULT resultid="1276" eventid="32" swimtime="00:01:15.43" lane="1" heatid="32002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1277" eventid="44" swimtime="00:00:31.41" lane="1" heatid="44002" />
                <RESULT resultid="1278" eventid="52" swimtime="00:02:49.76" lane="1" heatid="52001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                    <SPLIT distance="100" swimtime="00:01:23.11" />
                    <SPLIT distance="150" swimtime="00:02:08.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="281" birthdate="2008-01-01" gender="M" lastname="Selingr" firstname="Lukás" license="0">
              <RESULTS>
                <RESULT resultid="1279" eventid="30" swimtime="00:00:58.80" lane="2" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1280" eventid="32" swimtime="00:00:54.48" lane="2" heatid="32009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1281" eventid="42" swimtime="00:00:26.69" lane="2" heatid="42010" />
                <RESULT resultid="1282" eventid="44" swimtime="00:00:25.64" lane="1" heatid="44012" />
                <RESULT resultid="1283" eventid="50" swimtime="00:02:17.64" lane="2" heatid="50001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="100" swimtime="00:01:07.08" />
                    <SPLIT distance="150" swimtime="00:01:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1284" eventid="52" swimtime="00:01:59.22" lane="3" heatid="52005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="100" swimtime="00:00:58.64" />
                    <SPLIT distance="150" swimtime="00:01:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2086" eventid="66" swimtime="00:00:26.17" lane="4" heatid="66001" />
                <RESULT resultid="2099" eventid="69" swimtime="00:00:25.21" lane="4" heatid="69001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="282" birthdate="2006-01-01" gender="M" lastname="Werschall" firstname="Michal" license="0">
              <RESULTS>
                <RESULT resultid="1285" eventid="26" swimtime="00:00:28.98" lane="1" heatid="26010" />
                <RESULT resultid="1286" eventid="36" swimtime="00:02:21.61" lane="3" heatid="36002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1287" eventid="42" swimtime="00:00:29.07" lane="2" heatid="42006" />
                <RESULT resultid="1288" eventid="44" swimtime="00:00:27.05" lane="1" heatid="44008" />
                <RESULT resultid="1289" eventid="48" swimtime="00:01:03.88" lane="2" heatid="48005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2048" eventid="57" swimtime="00:00:28.41" lane="4" heatid="57001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="283" birthdate="2014-01-01" gender="F" lastname="Federselová" firstname="Ema" license="0">
              <RESULTS>
                <RESULT resultid="1290" eventid="3" swimtime="00:00:48.59" lane="4" heatid="3019" />
                <RESULT resultid="1291" eventid="7" swimtime="00:00:42.14" lane="4" heatid="7008" />
                <RESULT resultid="1292" eventid="15" swimtime="00:01:45.65" lane="4" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1293" eventid="19" swimtime="00:01:38.63" lane="3" heatid="19005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="284" birthdate="2014-01-01" gender="F" lastname="Kostolná" firstname="Alice" license="0">
              <RESULTS>
                <RESULT resultid="1294" eventid="3" swimtime="00:00:45.11" lane="2" heatid="3019" />
                <RESULT resultid="1295" eventid="9" swimtime="00:01:41.72" lane="2" heatid="9012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1296" eventid="15" swimtime="00:01:35.70" lane="2" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1297" eventid="19" swimtime="00:01:28.53" lane="3" heatid="19013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="285" birthdate="2014-01-01" gender="F" lastname="Meinlová" firstname="Tereza" license="0">
              <RESULTS>
                <RESULT resultid="1298" eventid="3" swimtime="00:00:43.83" lane="3" heatid="3019" />
                <RESULT resultid="1299" eventid="7" swimtime="00:00:41.58" lane="2" heatid="7010" />
                <RESULT resultid="1300" eventid="15" status="DSQ" swimtime="00:01:35.78" lane="3" heatid="15011" comment="Die Sportlerin hat bei der zweiten Wende nach Verlassen der Rückenlage nicht unverzüglich die eigentliche Wendenbewegung ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1301" eventid="19" swimtime="00:01:36.29" lane="3" heatid="19007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="286" birthdate="2014-01-01" gender="F" lastname="Ruzková" firstname="Ella" license="0">
              <RESULTS>
                <RESULT resultid="1302" eventid="7" swimtime="00:00:39.43" lane="2" heatid="7020" />
                <RESULT resultid="1303" eventid="9" swimtime="00:01:43.38" lane="3" heatid="9012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1304" eventid="13" swimtime="00:00:49.89" lane="3" heatid="13007" />
                <RESULT resultid="1305" eventid="19" swimtime="00:01:30.89" lane="2" heatid="19013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="287" birthdate="2012-01-01" gender="F" lastname="Dolezalová" firstname="Barbora" license="0">
              <RESULTS>
                <RESULT resultid="1306" eventid="3" swimtime="00:00:42.40" lane="3" heatid="3015" />
                <RESULT resultid="1307" eventid="5" swimtime="00:01:42.33" lane="4" heatid="5006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1308" eventid="7" swimtime="00:00:37.35" lane="1" heatid="7015" />
                <RESULT resultid="1309" eventid="15" swimtime="00:01:33.09" lane="3" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1310" eventid="17" swimtime="00:00:46.28" lane="3" heatid="17008" />
                <RESULT resultid="1311" eventid="19" swimtime="00:01:25.20" lane="1" heatid="19009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="288" birthdate="2012-01-01" gender="F" lastname="Hirsová" firstname="Nela" license="0">
              <RESULTS>
                <RESULT resultid="1312" eventid="3" status="DNS" swimtime="00:00:00.00" lane="3" heatid="3012" />
                <RESULT resultid="1313" eventid="5" status="DNS" swimtime="00:00:00.00" lane="4" heatid="5005" />
                <RESULT resultid="1314" eventid="7" status="DNS" swimtime="00:00:00.00" lane="3" heatid="7014" />
                <RESULT resultid="1315" eventid="13" status="DNS" swimtime="00:00:00.00" lane="4" heatid="13002" />
                <RESULT resultid="1316" eventid="17" status="DNS" swimtime="00:00:00.00" lane="4" heatid="17008" />
                <RESULT resultid="1317" eventid="19" status="DNS" swimtime="00:00:00.00" lane="2" heatid="19008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="289" birthdate="2012-01-01" gender="F" lastname="Jaklová" firstname="Valerie" license="0">
              <RESULTS>
                <RESULT resultid="1318" eventid="3" swimtime="00:00:39.09" lane="1" heatid="3021" />
                <RESULT resultid="1319" eventid="5" swimtime="00:01:54.15" lane="2" heatid="5004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1320" eventid="7" swimtime="00:00:35.35" lane="3" heatid="7017" />
                <RESULT resultid="1321" eventid="15" swimtime="00:01:26.11" lane="4" heatid="15013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1322" eventid="17" swimtime="00:00:52.69" lane="3" heatid="17006" />
                <RESULT resultid="1323" eventid="19" swimtime="00:01:17.35" lane="2" heatid="19010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="290" birthdate="2012-01-01" gender="F" lastname="Klánová" firstname="Stela" license="0">
              <RESULTS>
                <RESULT resultid="1324" eventid="1" status="DNS" swimtime="00:00:00.00" lane="2" heatid="1002" />
                <RESULT resultid="1325" eventid="3" swimtime="00:00:36.69" lane="2" heatid="3021" />
                <RESULT resultid="1326" eventid="7" swimtime="00:00:32.62" lane="2" heatid="7022" />
                <RESULT resultid="1327" eventid="13" swimtime="00:00:37.83" lane="4" heatid="13009" />
                <RESULT resultid="1328" eventid="15" swimtime="00:01:24.20" lane="1" heatid="15013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1329" eventid="19" swimtime="00:01:18.89" lane="2" heatid="19011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="291" birthdate="2012-01-01" gender="F" lastname="Kosatová" firstname="Veronika" license="0">
              <RESULTS>
                <RESULT resultid="1330" eventid="3" swimtime="00:00:37.46" lane="3" heatid="3021" />
                <RESULT resultid="1331" eventid="7" swimtime="00:00:33.75" lane="4" heatid="7022" />
                <RESULT resultid="1332" eventid="9" swimtime="00:01:24.61" lane="3" heatid="9014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1333" eventid="13" swimtime="00:00:40.50" lane="2" heatid="13005" />
                <RESULT resultid="1334" eventid="15" swimtime="00:01:23.04" lane="2" heatid="15013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1335" eventid="19" swimtime="00:01:15.01" lane="3" heatid="19015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="292" birthdate="2012-01-01" gender="F" lastname="Kvetová" firstname="Markéta" license="0">
              <RESULTS>
                <RESULT resultid="1336" eventid="3" swimtime="00:00:44.21" lane="2" heatid="3014" />
                <RESULT resultid="1337" eventid="7" swimtime="00:00:39.92" lane="2" heatid="7012" />
                <RESULT resultid="1338" eventid="9" swimtime="00:01:38.67" lane="2" heatid="9007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1339" eventid="13" swimtime="00:00:49.97" lane="1" heatid="13003" />
                <RESULT resultid="1340" eventid="15" swimtime="00:01:34.10" lane="4" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1341" eventid="19" swimtime="00:01:27.34" lane="1" heatid="19008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="293" birthdate="2012-01-01" gender="F" lastname="Legnerová" firstname="Jana" license="0">
              <RESULTS>
                <RESULT resultid="1342" eventid="3" swimtime="00:00:39.04" lane="2" heatid="3015" />
                <RESULT resultid="1343" eventid="7" swimtime="00:00:32.77" lane="3" heatid="7022" />
                <RESULT resultid="1344" eventid="9" swimtime="00:01:22.01" lane="2" heatid="9014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1345" eventid="13" swimtime="00:00:40.61" lane="4" heatid="13005" />
                <RESULT resultid="1346" eventid="19" swimtime="00:01:13.10" lane="2" heatid="19015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1347" eventid="21" swimtime="00:02:59.28" lane="2" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:01:26.88" />
                    <SPLIT distance="150" swimtime="00:02:19.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="294" birthdate="2012-01-01" gender="F" lastname="Steckerová" firstname="Klára" license="0">
              <RESULTS>
                <RESULT resultid="1348" eventid="3" swimtime="00:00:42.10" lane="2" heatid="3013" />
                <RESULT resultid="1349" eventid="5" swimtime="00:01:36.89" lane="1" heatid="5011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1350" eventid="7" swimtime="00:00:37.34" lane="1" heatid="7002" />
                <RESULT resultid="1351" eventid="13" swimtime="00:00:44.35" lane="1" heatid="13009" />
                <RESULT resultid="1352" eventid="17" swimtime="00:00:45.12" lane="4" heatid="17009" />
                <RESULT resultid="1353" eventid="19" swimtime="00:01:20.66" lane="1" heatid="19010">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="295" birthdate="2012-01-01" gender="F" lastname="Valesová" firstname="Josefína" license="0">
              <RESULTS>
                <RESULT resultid="1354" eventid="1" swimtime="00:01:39.35" lane="1" heatid="1001">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1355" eventid="5" swimtime="00:01:25.97" lane="2" heatid="5011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1356" eventid="9" swimtime="00:01:26.09" lane="4" heatid="9014">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1357" eventid="13" swimtime="00:00:41.16" lane="3" heatid="13005" />
                <RESULT resultid="1358" eventid="17" swimtime="00:00:39.56" lane="3" heatid="17013" />
                <RESULT resultid="1359" eventid="21" swimtime="00:03:08.98" lane="4" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:31.80" />
                    <SPLIT distance="150" swimtime="00:02:21.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="296" birthdate="2012-01-01" gender="F" lastname="Zaspalová" firstname="Nela" license="0">
              <RESULTS>
                <RESULT resultid="1360" eventid="3" swimtime="00:00:43.05" lane="4" heatid="3021" />
                <RESULT resultid="1361" eventid="5" swimtime="00:01:41.98" lane="2" heatid="5006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1362" eventid="7" swimtime="00:00:35.68" lane="4" heatid="7016" />
                <RESULT resultid="1363" eventid="15" swimtime="00:01:36.96" lane="1" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1364" eventid="17" swimtime="00:00:45.85" lane="4" heatid="17013" />
                <RESULT resultid="1365" eventid="19" swimtime="00:01:19.98" lane="2" heatid="19009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="297" birthdate="2011-01-01" gender="F" lastname="Tumová" firstname="Adéla" license="0">
              <RESULTS>
                <RESULT resultid="1366" eventid="3" swimtime="00:00:37.75" lane="2" heatid="3017" />
                <RESULT resultid="1367" eventid="7" swimtime="00:00:32.77" lane="3" heatid="7018" />
                <RESULT resultid="1368" eventid="9" swimtime="00:01:23.66" lane="3" heatid="9015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1369" eventid="15" swimtime="00:01:27.98" lane="2" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1370" eventid="17" swimtime="00:00:45.14" lane="1" heatid="17009" />
                <RESULT resultid="1371" eventid="19" swimtime="00:01:17.56" lane="1" heatid="19011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="298" birthdate="2013-01-01" gender="F" lastname="Sykorová" firstname="Zuzana" license="0">
              <RESULTS>
                <RESULT resultid="1372" eventid="3" swimtime="00:00:43.43" lane="4" heatid="3020" />
                <RESULT resultid="1373" eventid="7" swimtime="00:00:40.29" lane="4" heatid="7021" />
                <RESULT resultid="1374" eventid="9" swimtime="00:01:41.52" lane="4" heatid="9007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1375" eventid="15" swimtime="00:01:40.48" lane="3" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1376" eventid="17" swimtime="00:00:53.12" lane="4" heatid="17012" />
                <RESULT resultid="1377" eventid="19" swimtime="00:01:28.88" lane="3" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="299" birthdate="2015-01-01" gender="M" lastname="Dousa" firstname="Mikulás" license="0">
              <RESULTS>
                <RESULT resultid="1378" eventid="4" swimtime="00:00:40.52" lane="2" heatid="4010" />
                <RESULT resultid="1379" eventid="8" swimtime="00:00:35.52" lane="2" heatid="8015" />
                <RESULT resultid="1380" eventid="14" swimtime="00:00:48.69" lane="4" heatid="14003" />
                <RESULT resultid="1381" eventid="20" swimtime="00:01:23.40" lane="2" heatid="20011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="300" birthdate="2014-01-01" gender="M" lastname="Kundrát" firstname="Jan" license="0">
              <RESULTS>
                <RESULT resultid="1382" eventid="4" status="DNS" swimtime="00:00:00.00" lane="1" heatid="4011" />
                <RESULT resultid="1383" eventid="8" status="DNS" swimtime="00:00:00.00" lane="4" heatid="8016" />
                <RESULT resultid="1384" eventid="18" status="DNS" swimtime="00:00:00.00" lane="4" heatid="18009" />
                <RESULT resultid="1385" eventid="20" status="DNS" swimtime="00:00:00.00" lane="4" heatid="20012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="301" birthdate="2014-01-01" gender="M" lastname="Vales" firstname="Josef" license="0">
              <RESULTS>
                <RESULT resultid="1386" eventid="6" swimtime="00:01:39.61" lane="2" heatid="6006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1387" eventid="8" swimtime="00:00:34.07" lane="3" heatid="8016" />
                <RESULT resultid="1388" eventid="14" swimtime="00:00:38.19" lane="3" heatid="14007" />
                <RESULT resultid="1389" eventid="20" swimtime="00:01:18.05" lane="3" heatid="20012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="302" birthdate="2012-01-01" gender="M" lastname="Zák" firstname="Jiri" license="0">
              <RESULTS>
                <RESULT resultid="1390" eventid="4" swimtime="00:00:49.47" lane="1" heatid="4003" />
                <RESULT resultid="1391" eventid="8" swimtime="00:00:41.73" lane="1" heatid="8004" />
                <RESULT resultid="1392" eventid="16" status="DSQ" swimtime="00:01:46.25" lane="3" heatid="16002" comment="Der Sportler hat bei der ersten, zweiten und dritten Wende nach Verlassen der Rückenlage und Abschluss des Armzugs die eigentliche Wendenbewegung nicht unverzüglich ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1393" eventid="20" swimtime="00:01:38.82" lane="2" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="303" birthdate="2011-01-01" gender="M" lastname="Goncar" firstname="Daniel" license="0">
              <RESULTS>
                <RESULT resultid="1394" eventid="2" status="WDR" swimtime="00:00:00.00" lane="0" heatid="2000" />
                <RESULT resultid="1395" eventid="6" status="WDR" swimtime="00:00:00.00" lane="0" heatid="6000" />
                <RESULT resultid="1396" eventid="10" status="WDR" swimtime="00:00:00.00" lane="0" heatid="10000" />
                <RESULT resultid="1397" eventid="14" status="WDR" swimtime="00:00:00.00" lane="0" heatid="14000" />
                <RESULT resultid="1398" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="1399" eventid="18" status="WDR" swimtime="00:00:00.00" lane="0" heatid="18000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="304" birthdate="2011-01-01" gender="M" lastname="Hrych" firstname="Jan" license="0">
              <RESULTS>
                <RESULT resultid="1400" eventid="4" swimtime="00:00:43.26" lane="3" heatid="4008" />
                <RESULT resultid="1401" eventid="6" swimtime="00:01:48.67" lane="4" heatid="6009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1402" eventid="8" swimtime="00:00:37.87" lane="2" heatid="8010" />
                <RESULT resultid="1403" eventid="16" swimtime="00:01:35.40" lane="3" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1404" eventid="18" swimtime="00:00:49.90" lane="4" heatid="18006" />
                <RESULT resultid="1405" eventid="20" swimtime="00:01:27.34" lane="4" heatid="20015">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="305" birthdate="2011-01-01" gender="M" lastname="Vymetal" firstname="Oliver" license="0">
              <RESULTS>
                <RESULT resultid="1406" eventid="4" status="WDR" swimtime="00:00:00.00" lane="0" heatid="4000" />
                <RESULT resultid="1407" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="1408" eventid="10" status="WDR" swimtime="00:00:00.00" lane="0" heatid="10000" />
                <RESULT resultid="1409" eventid="14" status="WDR" swimtime="00:00:00.00" lane="0" heatid="14000" />
                <RESULT resultid="1410" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="1411" eventid="22" status="WDR" swimtime="00:00:00.00" lane="0" heatid="22000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="306" birthdate="2012-01-01" gender="M" lastname="Dousa" firstname="Matous" license="0">
              <RESULTS>
                <RESULT resultid="1412" eventid="4" swimtime="00:00:39.65" lane="1" heatid="4009" />
                <RESULT resultid="1413" eventid="6" swimtime="00:01:46.26" lane="1" heatid="6005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1414" eventid="8" swimtime="00:00:35.89" lane="1" heatid="8012" />
                <RESULT resultid="1415" eventid="16" swimtime="00:01:26.36" lane="4" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1416" eventid="18" swimtime="00:00:51.39" lane="3" heatid="18005" />
                <RESULT resultid="1417" eventid="20" swimtime="00:01:19.13" lane="2" heatid="20008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="307" birthdate="2012-01-01" gender="M" lastname="Masopust" firstname="Tomás" license="0">
              <RESULTS>
                <RESULT resultid="1418" eventid="2" status="WDR" swimtime="00:00:00.00" lane="0" heatid="2000" />
                <RESULT resultid="1419" eventid="6" status="WDR" swimtime="00:00:00.00" lane="0" heatid="6000" />
                <RESULT resultid="1420" eventid="8" status="WDR" swimtime="00:00:00.00" lane="0" heatid="8000" />
                <RESULT resultid="1421" eventid="14" status="WDR" swimtime="00:00:00.00" lane="0" heatid="14000" />
                <RESULT resultid="1422" eventid="16" status="WDR" swimtime="00:00:00.00" lane="0" heatid="16000" />
                <RESULT resultid="1423" eventid="18" status="WDR" swimtime="00:00:00.00" lane="0" heatid="18000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="308" birthdate="2012-01-01" gender="M" lastname="Krpálek" firstname="Tomás" license="0">
              <RESULTS>
                <RESULT resultid="1424" eventid="4" swimtime="00:00:46.14" lane="2" heatid="4005" />
                <RESULT resultid="1425" eventid="6" swimtime="00:01:59.30" lane="3" heatid="6003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1426" eventid="8" swimtime="00:00:38.63" lane="4" heatid="8012" />
                <RESULT resultid="1427" eventid="16" swimtime="00:01:43.62" lane="4" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1428" eventid="18" swimtime="00:00:52.95" lane="1" heatid="18005" />
                <RESULT resultid="1429" eventid="20" swimtime="00:01:32.41" lane="3" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="309" birthdate="2012-01-01" gender="M" lastname="Ziacek" firstname="Lukás" license="0">
              <RESULTS>
                <RESULT resultid="1430" eventid="4" swimtime="00:00:45.06" lane="3" heatid="4006" />
                <RESULT resultid="1431" eventid="6" swimtime="00:01:54.20" lane="2" heatid="6003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1432" eventid="8" swimtime="00:00:41.12" lane="2" heatid="8009" />
                <RESULT resultid="1433" eventid="16" swimtime="00:01:38.64" lane="1" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1434" eventid="18" swimtime="00:00:52.43" lane="2" heatid="18003" />
                <RESULT resultid="1435" eventid="20" swimtime="00:01:27.85" lane="4" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="310" birthdate="2013-01-01" gender="M" lastname="Kopta" firstname="Filip" license="0">
              <RESULTS>
                <RESULT resultid="1436" eventid="4" swimtime="00:00:41.02" lane="1" heatid="4012" />
                <RESULT resultid="1437" eventid="6" swimtime="00:01:47.73" lane="3" heatid="6005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1438" eventid="8" swimtime="00:00:37.15" lane="2" heatid="8011" />
                <RESULT resultid="1439" eventid="16" swimtime="00:01:31.77" lane="4" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1440" eventid="18" swimtime="00:00:49.70" lane="4" heatid="18010" />
                <RESULT resultid="1441" eventid="20" swimtime="00:01:23.62" lane="4" heatid="20008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="311" birthdate="2013-01-01" gender="M" lastname="Krecek" firstname="Jáchym" license="0">
              <RESULTS>
                <RESULT resultid="1442" eventid="2" swimtime="00:01:28.51" lane="2" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1443" eventid="8" swimtime="00:00:35.21" lane="3" heatid="8017" />
                <RESULT resultid="1444" eventid="10" swimtime="00:01:29.56" lane="3" heatid="10008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1445" eventid="14" swimtime="00:00:37.07" lane="2" heatid="14008" />
                <RESULT resultid="1446" eventid="16" swimtime="00:01:28.43" lane="2" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1447" eventid="20" swimtime="00:01:18.78" lane="1" heatid="20013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="312" birthdate="2013-01-01" gender="M" lastname="Kyncl" firstname="Ondrej" license="0">
              <RESULTS>
                <RESULT resultid="1448" eventid="2" swimtime="00:01:36.13" lane="3" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1449" eventid="4" status="DSQ" swimtime="00:00:38.32" lane="2" heatid="4012" comment="Der Sportler startete vor dem Startsignal" />
                <RESULT resultid="1450" eventid="8" swimtime="00:00:34.39" lane="2" heatid="8017" />
                <RESULT resultid="1451" eventid="14" swimtime="00:00:38.17" lane="1" heatid="14008" />
                <RESULT resultid="1452" eventid="16" swimtime="00:01:23.42" lane="3" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1453" eventid="20" swimtime="00:01:14.69" lane="2" heatid="20013">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="313" birthdate="2013-01-01" gender="M" lastname="Rybár" firstname="Vojtech" license="0">
              <RESULTS>
                <RESULT resultid="1454" eventid="2" swimtime="00:01:30.92" lane="1" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1455" eventid="6" swimtime="00:01:39.50" lane="1" heatid="6007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1456" eventid="10" swimtime="00:01:25.49" lane="2" heatid="10008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1457" eventid="14" swimtime="00:00:38.82" lane="3" heatid="14008" />
                <RESULT resultid="1458" eventid="20" status="DNS" swimtime="00:00:00.00" lane="3" heatid="20013" />
                <RESULT resultid="1459" eventid="22" status="DNS" swimtime="00:00:00.00" lane="3" heatid="22002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="314" birthdate="2013-01-01" gender="M" lastname="Weinhofer" firstname="Petr" license="0">
              <RESULTS>
                <RESULT resultid="1460" eventid="4" status="DNS" swimtime="00:00:00.00" lane="1" heatid="4007" />
                <RESULT resultid="1461" eventid="6" status="DNS" swimtime="00:00:00.00" lane="2" heatid="6004" />
                <RESULT resultid="1462" eventid="8" status="DNS" swimtime="00:00:00.00" lane="3" heatid="8012" />
                <RESULT resultid="1463" eventid="14" status="DNS" swimtime="00:00:00.00" lane="1" heatid="14002" />
                <RESULT resultid="1464" eventid="18" status="DNS" swimtime="00:00:00.00" lane="1" heatid="18010" />
                <RESULT resultid="1465" eventid="20" status="DNS" swimtime="00:00:00.00" lane="1" heatid="20007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="414" birthdate="2009-01-01" gender="M" lastname="Pechác" firstname="Denis" license="0">
              <RESULTS>
                <RESULT resultid="1940" eventid="26" swimtime="00:00:34.70" lane="4" heatid="26008" />
                <RESULT resultid="1941" eventid="32" swimtime="00:01:07.86" lane="4" heatid="32008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1942" eventid="34" swimtime="00:01:17.99" lane="1" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1943" eventid="42" swimtime="00:00:35.88" lane="2" heatid="42001" />
                <RESULT resultid="1944" eventid="44" swimtime="00:00:30.39" lane="3" heatid="44002" />
                <RESULT resultid="1945" eventid="48" swimtime="00:01:14.29" lane="2" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1466" eventid="11" swimtime="00:02:18.50" lane="3" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:06.88" />
                    <SPLIT distance="150" swimtime="00:01:41.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="289" number="1" />
                    <RELAYPOSITION athleteid="293" number="2" />
                    <RELAYPOSITION athleteid="301" number="3" />
                    <RELAYPOSITION athleteid="309" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1467" eventid="23" swimtime="00:02:37.92" lane="4" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:21.56" />
                    <SPLIT distance="150" swimtime="00:01:58.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="306" number="1" />
                    <RELAYPOSITION athleteid="295" number="2" />
                    <RELAYPOSITION athleteid="290" number="3" />
                    <RELAYPOSITION athleteid="308" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1468" eventid="11" swimtime="00:02:18.80" lane="1" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:43.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="299" number="1" />
                    <RELAYPOSITION athleteid="291" number="2" />
                    <RELAYPOSITION athleteid="296" number="3" />
                    <RELAYPOSITION athleteid="304" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1469" eventid="23" swimtime="00:03:00.35" lane="1" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                    <SPLIT distance="100" swimtime="00:01:29.83" />
                    <SPLIT distance="150" swimtime="00:02:20.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="284" number="1" />
                    <RELAYPOSITION athleteid="301" number="2" />
                    <RELAYPOSITION athleteid="286" number="3" />
                    <RELAYPOSITION athleteid="302" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1470" eventid="39" swimtime="00:01:56.34" lane="1" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:00:59.18" />
                    <SPLIT distance="150" swimtime="00:01:27.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="271" number="1" />
                    <RELAYPOSITION athleteid="272" number="2" />
                    <RELAYPOSITION athleteid="273" number="3" />
                    <RELAYPOSITION athleteid="266" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1471" eventid="71" swimtime="00:02:05.14" lane="1" heatid="71001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:36.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="266" number="1" />
                    <RELAYPOSITION athleteid="271" number="2" />
                    <RELAYPOSITION athleteid="273" number="3" />
                    <RELAYPOSITION athleteid="272" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1472" eventid="39" status="DNS" swimtime="00:00:00.00" lane="3" heatid="39001" />
                <RESULT resultid="1473" eventid="71" status="DNS" swimtime="00:00:00.00" lane="3" heatid="71001" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1474" eventid="40" swimtime="00:01:43.83" lane="3" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.90" />
                    <SPLIT distance="100" swimtime="00:00:51.37" />
                    <SPLIT distance="150" swimtime="00:01:17.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="278" number="1" />
                    <RELAYPOSITION athleteid="279" number="2" />
                    <RELAYPOSITION athleteid="282" number="3" />
                    <RELAYPOSITION athleteid="281" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1475" eventid="72" swimtime="00:01:50.45" lane="3" heatid="72001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                    <SPLIT distance="100" swimtime="00:00:58.91" />
                    <SPLIT distance="150" swimtime="00:01:25.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="282" number="1" />
                    <RELAYPOSITION athleteid="279" number="2" />
                    <RELAYPOSITION athleteid="281" number="3" />
                    <RELAYPOSITION athleteid="278" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1476" eventid="40" swimtime="00:01:54.77" lane="2" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="100" swimtime="00:00:57.23" />
                    <SPLIT distance="150" swimtime="00:01:26.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="277" number="1" />
                    <RELAYPOSITION athleteid="280" number="2" />
                    <RELAYPOSITION athleteid="414" number="3" />
                    <RELAYPOSITION athleteid="276" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1477" eventid="72" swimtime="00:02:06.44" lane="1" heatid="72001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="100" swimtime="00:01:01.95" />
                    <SPLIT distance="150" swimtime="00:01:35.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="277" number="1" />
                    <RELAYPOSITION athleteid="276" number="2" />
                    <RELAYPOSITION athleteid="414" number="3" />
                    <RELAYPOSITION athleteid="280" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TJ Slavie VS Plzen" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="323" birthdate="2006-01-01" gender="F" lastname="Studentová" firstname="Valentýna" license="0">
              <RESULTS>
                <RESULT resultid="1485" eventid="27" status="WDR" swimtime="00:00:00.00" lane="0" heatid="27000" />
                <RESULT resultid="1486" eventid="37" status="WDR" swimtime="00:00:00.00" lane="0" heatid="37000" />
                <RESULT resultid="1487" eventid="45" status="WDR" swimtime="00:00:00.00" lane="0" heatid="45000" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSV Einheit Süd Chemnitz e.V." nation="GER" region="12" code="3403">
          <ATHLETES>
            <ATHLETE athleteid="236" birthdate="2008-01-01" gender="F" lastname="Brabenetz" firstname="Jenna" license="393444">
              <RESULTS>
                <RESULT resultid="1105" eventid="25" swimtime="00:00:40.69" lane="1" heatid="25003" />
                <RESULT resultid="1106" eventid="29" swimtime="00:01:29.86" lane="3" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1107" eventid="31" swimtime="00:01:20.58" lane="3" heatid="31002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1108" eventid="43" swimtime="00:00:35.52" lane="3" heatid="43003" />
                <RESULT resultid="1109" eventid="47" swimtime="00:01:31.73" lane="1" heatid="47003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="237" birthdate="2008-01-01" gender="F" lastname="Hänig" firstname="Lilly" license="428120">
              <RESULTS>
                <RESULT resultid="1110" eventid="27" status="DSQ" swimtime="00:00:43.05" lane="2" heatid="27002" comment="Nach der Wende hat die Sportlerin mehrere Beinschläge ausgeführt." />
                <RESULT resultid="1111" eventid="31" swimtime="00:01:21.62" lane="4" heatid="31004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1112" eventid="37" swimtime="00:03:38.61" lane="4" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="100" swimtime="00:01:44.08" />
                    <SPLIT distance="150" swimtime="00:02:41.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1113" eventid="45" swimtime="00:01:38.06" lane="1" heatid="45001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="238" birthdate="2006-01-01" gender="F" lastname="Köhler" firstname="Lea Sophie" license="387692">
              <RESULTS>
                <RESULT resultid="1114" eventid="29" swimtime="00:01:15.76" lane="2" heatid="29006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1115" eventid="31" swimtime="00:01:06.71" lane="3" heatid="31012">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1116" eventid="41" swimtime="00:00:32.08" lane="4" heatid="41013" />
                <RESULT resultid="1117" eventid="43" swimtime="00:00:30.11" lane="4" heatid="43016" />
                <RESULT resultid="1118" eventid="47" swimtime="00:01:22.16" lane="3" heatid="47009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="239" birthdate="1992-01-01" gender="M" lastname="Metzner" firstname="Joshua" license="149240">
              <RESULTS>
                <RESULT resultid="1119" eventid="26" swimtime="00:00:29.71" lane="4" heatid="26007" />
                <RESULT resultid="1120" eventid="54" swimtime="00:02:21.95" lane="3" heatid="54003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                    <SPLIT distance="100" swimtime="00:01:06.94" />
                    <SPLIT distance="150" swimtime="00:01:48.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="240" birthdate="2009-01-01" gender="F" lastname="Rudolph" firstname="Anna" license="386529">
              <RESULTS>
                <RESULT resultid="1121" eventid="27" swimtime="00:00:43.94" lane="3" heatid="27002" />
                <RESULT resultid="1122" eventid="31" swimtime="00:01:23.09" lane="2" heatid="31002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1123" eventid="41" swimtime="00:00:42.72" lane="1" heatid="41001" />
                <RESULT resultid="1124" eventid="43" swimtime="00:00:36.84" lane="1" heatid="43003" />
                <RESULT resultid="1125" eventid="51" swimtime="00:03:06.91" lane="1" heatid="51002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:01:28.73" />
                    <SPLIT distance="150" swimtime="00:02:19.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="241" birthdate="2008-01-01" gender="F" lastname="Süß" firstname="Julia" license="391096">
              <RESULTS>
                <RESULT resultid="1126" eventid="25" swimtime="00:00:41.00" lane="1" heatid="25002" />
                <RESULT resultid="1127" eventid="29" swimtime="00:01:26.88" lane="2" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1128" eventid="31" swimtime="00:01:16.77" lane="1" heatid="31004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1129" eventid="41" swimtime="00:00:36.98" lane="4" heatid="41004" />
                <RESULT resultid="1130" eventid="43" swimtime="00:00:35.07" lane="3" heatid="43005" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Ústecká akademie plaveckých sportu" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="258" birthdate="2004-01-01" gender="M" lastname="Beca" firstname="Jakub" license="0">
              <RESULTS>
                <RESULT resultid="1170" eventid="26" swimtime="00:00:27.33" lane="3" heatid="26011" />
                <RESULT resultid="1171" eventid="32" swimtime="00:00:54.34" lane="2" heatid="32011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1172" eventid="36" swimtime="00:02:16.48" lane="2" heatid="36002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:42.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1173" eventid="42" swimtime="00:00:26.26" lane="1" heatid="42012" />
                <RESULT resultid="1174" eventid="44" swimtime="00:00:24.42" lane="1" heatid="44014" />
                <RESULT resultid="1175" eventid="48" swimtime="00:00:59.60" lane="3" heatid="48006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2050" eventid="58" swimtime="00:00:26.91" lane="3" heatid="58001" />
                <RESULT resultid="2085" eventid="66" swimtime="00:00:25.89" lane="1" heatid="66001" />
                <RESULT resultid="2103" eventid="70" swimtime="00:00:24.17" lane="4" heatid="70001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="259" birthdate="2008-01-01" gender="M" lastname="Bartuska" firstname="Daniel" license="0">
              <RESULTS>
                <RESULT resultid="1176" eventid="32" swimtime="00:01:01.48" lane="1" heatid="32006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1177" eventid="38" swimtime="00:02:47.22" lane="4" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:05.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1178" eventid="42" swimtime="00:00:30.19" lane="4" heatid="42010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="260" birthdate="2008-01-01" gender="F" lastname="Boriková" firstname="Barbora" license="0">
              <RESULTS>
                <RESULT resultid="1179" eventid="25" swimtime="00:00:33.21" lane="3" heatid="25008" />
                <RESULT resultid="1180" eventid="27" swimtime="00:00:36.77" lane="3" heatid="27007" />
                <RESULT resultid="1181" eventid="43" swimtime="00:00:30.03" lane="1" heatid="43015" />
                <RESULT resultid="1182" eventid="45" swimtime="00:01:20.78" lane="2" heatid="45005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2053" eventid="59" swimtime="00:00:36.69" lane="2" heatid="59001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="261" birthdate="2008-01-01" gender="F" lastname="Krivánková" firstname="Veronika" license="0">
              <RESULTS>
                <RESULT resultid="1183" eventid="25" swimtime="00:00:38.53" lane="3" heatid="25004" />
                <RESULT resultid="1184" eventid="27" swimtime="00:00:39.90" lane="1" heatid="27007" />
                <RESULT resultid="1185" eventid="37" swimtime="00:02:55.84" lane="2" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:24.51" />
                    <SPLIT distance="150" swimtime="00:02:10.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1186" eventid="43" swimtime="00:00:32.57" lane="4" heatid="43007" />
                <RESULT resultid="1187" eventid="45" swimtime="00:01:24.41" lane="3" heatid="45005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1188" eventid="47" swimtime="00:01:24.03" lane="1" heatid="47005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="262" birthdate="2008-01-01" gender="F" lastname="Gaberová" firstname="Alzbeta" license="0">
              <RESULTS>
                <RESULT resultid="1189" eventid="25" swimtime="00:00:35.06" lane="4" heatid="25007" />
                <RESULT resultid="1190" eventid="31" swimtime="00:01:06.76" lane="4" heatid="31008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1191" eventid="35" swimtime="00:02:34.75" lane="4" heatid="35003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:54.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1192" eventid="43" swimtime="00:00:31.01" lane="2" heatid="43007" />
                <RESULT resultid="1193" eventid="47" swimtime="00:01:13.96" lane="4" heatid="47008">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="263" birthdate="2008-01-01" gender="F" lastname="Fleková" firstname="Marie" license="0">
              <RESULTS>
                <RESULT resultid="1194" eventid="27" status="DSQ" swimtime="00:00:38.85" lane="4" heatid="27007" comment="Nach dem Start hat die Sportlerin zwei Delphinbeinschläge ausgeführt." />
                <RESULT resultid="1195" eventid="31" swimtime="00:01:11.75" lane="3" heatid="31006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1196" eventid="37" swimtime="00:03:04.36" lane="3" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:27.53" />
                    <SPLIT distance="150" swimtime="00:02:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1197" eventid="45" swimtime="00:01:23.94" lane="4" heatid="45005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="264" birthdate="2008-01-01" gender="F" lastname="Salounová" firstname="Gábina" license="0">
              <RESULTS>
                <RESULT resultid="1198" eventid="29" swimtime="00:01:14.19" lane="2" heatid="29002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1199" eventid="37" swimtime="00:03:00.42" lane="1" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:26.51" />
                    <SPLIT distance="150" swimtime="00:02:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1200" eventid="45" swimtime="00:01:24.27" lane="1" heatid="45005">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1201" eventid="49" swimtime="00:02:48.17" lane="4" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:19.34" />
                    <SPLIT distance="150" swimtime="00:02:04.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="265" birthdate="2001-01-01" gender="M" lastname="Grupác" firstname="Radek" license="0">
              <RESULTS>
                <RESULT resultid="1202" eventid="28" swimtime="00:00:29.77" lane="4" heatid="28001" />
                <RESULT resultid="2066" eventid="62" status="WDR" swimtime="00:00:00.00" lane="0" heatid="62000" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="WSG Jena-Lobeda e.V." nation="GER" region="16" code="3278">
          <ATHLETES>
            <ATHLETE athleteid="5" birthdate="2010-01-01" gender="F" lastname="Grimmer" firstname="Rita" license="446916">
              <RESULTS>
                <RESULT resultid="26" eventid="31" swimtime="00:01:19.02" lane="4" heatid="31009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="27" eventid="33" swimtime="00:01:37.88" lane="4" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="28" eventid="43" swimtime="00:00:35.16" lane="4" heatid="43003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="6" birthdate="2010-01-01" gender="F" lastname="Klemm" firstname="Zoè Amelie" license="423552">
              <RESULTS>
                <RESULT resultid="29" eventid="27" swimtime="00:00:41.37" lane="2" heatid="27005" />
                <RESULT resultid="30" eventid="33" swimtime="00:01:26.82" lane="4" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="31" eventid="45" swimtime="00:01:34.15" lane="2" heatid="45003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="7" birthdate="2010-01-01" gender="M" lastname="Kovezin" firstname="Vladimir" license="423550">
              <RESULTS>
                <RESULT resultid="32" eventid="4" swimtime="00:00:39.02" lane="3" heatid="4009" />
                <RESULT resultid="33" eventid="8" swimtime="00:00:31.35" lane="4" heatid="8014" />
                <RESULT resultid="34" eventid="22" swimtime="00:03:14.84" lane="4" heatid="22003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                    <SPLIT distance="100" swimtime="00:01:32.89" />
                    <SPLIT distance="150" swimtime="00:02:31.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="8" birthdate="2011-01-01" gender="F" lastname="Mutschke" firstname="Luisa" license="442362">
              <RESULTS>
                <RESULT resultid="35" eventid="3" swimtime="00:00:42.25" lane="4" heatid="3015" />
                <RESULT resultid="36" eventid="9" swimtime="00:01:34.46" lane="1" heatid="9009">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="37" eventid="13" swimtime="00:00:45.44" lane="1" heatid="13004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="9" birthdate="2009-01-01" gender="M" lastname="Neuhaus" firstname="Jakob Friedrich" license="437045">
              <RESULTS>
                <RESULT resultid="38" eventid="26" swimtime="00:00:38.72" lane="1" heatid="26002" />
                <RESULT resultid="39" eventid="34" swimtime="00:01:24.87" lane="3" heatid="34001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="40" eventid="54" swimtime="00:03:05.64" lane="1" heatid="54001">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:26.71" />
                    <SPLIT distance="150" swimtime="00:02:24.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="10" birthdate="2010-01-01" gender="F" lastname="Schirmer" firstname="Pauline" license="423553">
              <RESULTS>
                <RESULT resultid="41" eventid="29" swimtime="00:01:48.34" lane="4" heatid="29003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="42" eventid="33" swimtime="00:01:30.67" lane="1" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="43" eventid="47" swimtime="00:01:29.01" lane="4" heatid="47006">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="11" birthdate="2011-01-01" gender="M" lastname="Simon" firstname="Bruno" license="442369">
              <RESULTS>
                <RESULT resultid="44" eventid="4" status="DNS" swimtime="00:00:00.00" lane="4" heatid="4014" />
                <RESULT resultid="45" eventid="10" status="DNS" swimtime="00:00:00.00" lane="3" heatid="10002" />
                <RESULT resultid="46" eventid="14" status="DNS" swimtime="00:00:00.00" lane="3" heatid="14002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="12" birthdate="2002-01-01" gender="M" lastname="Spörl" firstname="Nils" license="310433">
              <RESULTS>
                <RESULT resultid="47" eventid="32" swimtime="00:01:00.44" lane="4" heatid="32011">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="48" eventid="48" swimtime="00:01:08.78" lane="3" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="13" birthdate="2011-01-01" gender="F" lastname="Steiniger" firstname="Enne Therese" license="442367">
              <RESULTS>
                <RESULT resultid="49" eventid="3" swimtime="00:00:43.24" lane="4" heatid="3017" />
                <RESULT resultid="50" eventid="7" swimtime="00:00:35.09" lane="1" heatid="7016" />
                <RESULT resultid="51" eventid="21" swimtime="00:03:30.57" lane="1" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:37.75" />
                    <SPLIT distance="150" swimtime="00:02:43.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
